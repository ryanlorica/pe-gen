module MulAddRecFNToRaw_preMul(
    input [1:0] io_op,
    input [64:0] io_a,
    input [64:0] io_b,
    input [64:0] io_c,
    output[52:0] io_mulAddA,
    output[52:0] io_mulAddB,
    output[105:0] io_mulAddC,
    output io_toPostMul_isSigNaNAny,
    output io_toPostMul_isNaNAOrB,
    output io_toPostMul_isInfA,
    output io_toPostMul_isZeroA,
    output io_toPostMul_isInfB,
    output io_toPostMul_isZeroB,
    output io_toPostMul_signProd,
    output io_toPostMul_isNaNC,
    output io_toPostMul_isInfC,
    output io_toPostMul_isZeroC,
    output[12:0] io_toPostMul_sExpSum,
    output io_toPostMul_doSubMags,
    output io_toPostMul_CIsDominant,
    output[5:0] io_toPostMul_CDom_CAlignDist,
    output[54:0] io_toPostMul_highAlignedSigC,
    output io_toPostMul_bit0AlignedSigC
);

  wire T0;
  wire[162:0] alignedSigC;
  wire T1;
  wire T2;
  wire reduced4CExtra;
  wire[13:0] T3;
  wire[13:0] T190;
  wire[12:0] T4;
  wire[4:0] T5;
  wire T6;
  wire[4:0] T7;
  wire[12:0] T8;
  wire[64:0] T9;
  wire[5:0] T10;
  wire[7:0] CAlignDist;
  wire[7:0] T11;
  wire[7:0] T12;
  wire[12:0] posNatCAlignDist;
  wire[14:0] sNatCAlignDist;
  wire[13:0] T191;
  wire[12:0] rawC_sExp;
  wire[12:0] T13;
  wire[12:0] T14;
  wire[11:0] T15;
  wire T192;
  wire[14:0] sExpAlignedProd;
  wire[14:0] T16;
  wire[13:0] T193;
  wire[12:0] rawB_sExp;
  wire[12:0] T17;
  wire[12:0] T18;
  wire[11:0] T19;
  wire T194;
  wire[13:0] T195;
  wire[12:0] rawA_sExp;
  wire[12:0] T20;
  wire[12:0] T21;
  wire[11:0] T22;
  wire T196;
  wire T23;
  wire isMinCAlign;
  wire T24;
  wire T25;
  wire rawB_isZero;
  wire T26;
  wire[2:0] T27;
  wire rawA_isZero;
  wire T28;
  wire[2:0] T29;
  wire[3:0] T30;
  wire[1:0] T31;
  wire T32;
  wire[1:0] T33;
  wire[3:0] T34;
  wire T35;
  wire[1:0] T36;
  wire T37;
  wire[1:0] T38;
  wire T39;
  wire[7:0] T40;
  wire[7:0] T41;
  wire[7:0] T42;
  wire[6:0] T43;
  wire[7:0] T44;
  wire[7:0] T45;
  wire[7:0] T46;
  wire[5:0] T47;
  wire[7:0] T48;
  wire[7:0] T49;
  wire[7:0] T50;
  wire[3:0] T51;
  wire[7:0] T52;
  wire[7:0] T53;
  wire[7:0] T197;
  wire[3:0] T54;
  wire[7:0] T55;
  wire[7:0] T198;
  wire[5:0] T56;
  wire[7:0] T57;
  wire[7:0] T199;
  wire[6:0] T58;
  wire[13:0] T59;
  wire[13:0] T60;
  wire[6:0] T61;
  wire[3:0] T62;
  wire[1:0] T63;
  wire T64;
  wire T65;
  wire[3:0] T66;
  wire[53:0] T67;
  wire[53:0] rawC_sig;
  wire[53:0] T68;
  wire[52:0] T69;
  wire[51:0] T70;
  wire T71;
  wire T72;
  wire[2:0] T73;
  wire T74;
  wire T75;
  wire[3:0] T76;
  wire[1:0] T77;
  wire T78;
  wire T79;
  wire[3:0] T80;
  wire T81;
  wire T82;
  wire[3:0] T83;
  wire[2:0] T84;
  wire[1:0] T85;
  wire T86;
  wire T87;
  wire[3:0] T88;
  wire T89;
  wire T90;
  wire[3:0] T91;
  wire T92;
  wire T93;
  wire[3:0] T94;
  wire[6:0] T95;
  wire[3:0] T96;
  wire[1:0] T97;
  wire T98;
  wire T99;
  wire[3:0] T100;
  wire T101;
  wire T102;
  wire[3:0] T103;
  wire[1:0] T104;
  wire T105;
  wire T106;
  wire[3:0] T107;
  wire T108;
  wire T109;
  wire[3:0] T110;
  wire[2:0] T111;
  wire[1:0] T112;
  wire T113;
  wire T114;
  wire[3:0] T115;
  wire T116;
  wire T117;
  wire[3:0] T118;
  wire T119;
  wire T120;
  wire[1:0] T121;
  wire T122;
  wire[2:0] T123;
  wire[164:0] mainAlignedSigC;
  wire[164:0] T124;
  wire[164:0] T125;
  wire[110:0] T126;
  wire[110:0] T200;
  wire[53:0] T127;
  wire[53:0] T128;
  wire T129;
  wire T130;
  wire T131;
  wire[2:0] T132;
  wire doSubMags;
  wire T133;
  wire T134;
  wire rawC_sign;
  wire T135;
  wire signProd;
  wire T136;
  wire T137;
  wire rawB_sign;
  wire T138;
  wire rawA_sign;
  wire T139;
  wire[161:0] T140;
  wire[54:0] T141;
  wire[5:0] T142;
  wire CIsDominant;
  wire T143;
  wire T144;
  wire T145;
  wire rawC_isZero;
  wire[12:0] T201;
  wire[14:0] T146;
  wire[14:0] T147;
  wire[13:0] T202;
  wire T203;
  wire rawC_isInf;
  wire T148;
  wire T149;
  wire T150;
  wire T151;
  wire[1:0] T152;
  wire rawC_isNaN;
  wire T153;
  wire T154;
  wire rawB_isInf;
  wire T155;
  wire T156;
  wire T157;
  wire T158;
  wire[1:0] T159;
  wire rawA_isInf;
  wire T160;
  wire T161;
  wire T162;
  wire T163;
  wire[1:0] T164;
  wire T165;
  wire rawB_isNaN;
  wire T166;
  wire T167;
  wire rawA_isNaN;
  wire T168;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire T173;
  wire T174;
  wire T175;
  wire T176;
  wire T177;
  wire[53:0] rawB_sig;
  wire[53:0] T178;
  wire[52:0] T179;
  wire[51:0] T180;
  wire T181;
  wire T182;
  wire T183;
  wire T184;
  wire[53:0] rawA_sig;
  wire[53:0] T185;
  wire[52:0] T186;
  wire[51:0] T187;
  wire T188;
  wire[105:0] T189;
  wire[52:0] T204;
  wire[52:0] T205;


  assign io_toPostMul_bit0AlignedSigC = T0;
  assign T0 = alignedSigC[0];
  assign alignedSigC = {T140, T1};
  assign T1 = doSubMags ? T129 : T2;
  assign T2 = T122 | reduced4CExtra;
  assign reduced4CExtra = T3 != 14'h0;
  assign T3 = T59 & T190;
  assign T190 = {1'h0, T4};
  assign T4 = {T40, T5};
  assign T5 = {T30, T6};
  assign T6 = T7[4];
  assign T7 = T8[12:8];
  assign T8 = T9[36:24];
  assign T9 = $signed(65'h10000000000000000) >>> T10;
  assign T10 = CAlignDist >> 2'h2;
  assign CAlignDist = isMinCAlign ? 8'h0 : T11;
  assign T11 = T23 ? T12 : 8'ha1;
  assign T12 = posNatCAlignDist[7:0];
  assign posNatCAlignDist = sNatCAlignDist[12:0];
  assign sNatCAlignDist = sExpAlignedProd - T191;
  assign T191 = {T192, rawC_sExp};
  assign rawC_sExp = T13;
  assign T13 = T14;
  assign T14 = {1'h0, T15};
  assign T15 = io_c[63:52];
  assign T192 = rawC_sExp[12];
  assign sExpAlignedProd = T16 + 14'h3838;
  assign T16 = T195 + T193;
  assign T193 = {T194, rawB_sExp};
  assign rawB_sExp = T17;
  assign T17 = T18;
  assign T18 = {1'h0, T19};
  assign T19 = io_b[63:52];
  assign T194 = rawB_sExp[12];
  assign T195 = {T196, rawA_sExp};
  assign rawA_sExp = T20;
  assign T20 = T21;
  assign T21 = {1'h0, T22};
  assign T22 = io_a[63:52];
  assign T196 = rawA_sExp[12];
  assign T23 = posNatCAlignDist < 13'ha1;
  assign isMinCAlign = T25 | T24;
  assign T24 = $signed(sNatCAlignDist) < $signed(1'h0);
  assign T25 = rawA_isZero | rawB_isZero;
  assign rawB_isZero = T26;
  assign T26 = T27 == 3'h0;
  assign T27 = T19[11:9];
  assign rawA_isZero = T28;
  assign T28 = T29 == 3'h0;
  assign T29 = T22[11:9];
  assign T30 = {T36, T31};
  assign T31 = {T35, T32};
  assign T32 = T33[1];
  assign T33 = T34[3:2];
  assign T34 = T7[3:0];
  assign T35 = T33[0];
  assign T36 = {T39, T37};
  assign T37 = T38[1];
  assign T38 = T34[1:0];
  assign T39 = T38[0];
  assign T40 = T57 | T41;
  assign T41 = T42 & 8'haa;
  assign T42 = T43 << 1'h1;
  assign T43 = T44[6:0];
  assign T44 = T55 | T45;
  assign T45 = T46 & 8'hcc;
  assign T46 = T47 << 2'h2;
  assign T47 = T48[5:0];
  assign T48 = T53 | T49;
  assign T49 = T50 & 8'hf0;
  assign T50 = T51 << 3'h4;
  assign T51 = T52[3:0];
  assign T52 = T8[7:0];
  assign T53 = T197 & 8'hf;
  assign T197 = {4'h0, T54};
  assign T54 = T52 >> 3'h4;
  assign T55 = T198 & 8'h33;
  assign T198 = {2'h0, T56};
  assign T56 = T48 >> 2'h2;
  assign T57 = T199 & 8'h55;
  assign T199 = {1'h0, T58};
  assign T58 = T44 >> 1'h1;
  assign T59 = T60;
  assign T60 = {T95, T61};
  assign T61 = {T84, T62};
  assign T62 = {T77, T63};
  assign T63 = {T74, T64};
  assign T64 = T65;
  assign T65 = T66 != 4'h0;
  assign T66 = T67[3:0];
  assign T67 = rawC_sig << 1'h0;
  assign rawC_sig = T68;
  assign T68 = {1'h0, T69};
  assign T69 = {T71, T70};
  assign T70 = io_c[51:0];
  assign T71 = T72 ^ 1'h1;
  assign T72 = T73 == 3'h0;
  assign T73 = T15[11:9];
  assign T74 = T75;
  assign T75 = T76 != 4'h0;
  assign T76 = T67[7:4];
  assign T77 = {T81, T78};
  assign T78 = T79;
  assign T79 = T80 != 4'h0;
  assign T80 = T67[11:8];
  assign T81 = T82;
  assign T82 = T83 != 4'h0;
  assign T83 = T67[15:12];
  assign T84 = {T92, T85};
  assign T85 = {T89, T86};
  assign T86 = T87;
  assign T87 = T88 != 4'h0;
  assign T88 = T67[19:16];
  assign T89 = T90;
  assign T90 = T91 != 4'h0;
  assign T91 = T67[23:20];
  assign T92 = T93;
  assign T93 = T94 != 4'h0;
  assign T94 = T67[27:24];
  assign T95 = {T111, T96};
  assign T96 = {T104, T97};
  assign T97 = {T101, T98};
  assign T98 = T99;
  assign T99 = T100 != 4'h0;
  assign T100 = T67[31:28];
  assign T101 = T102;
  assign T102 = T103 != 4'h0;
  assign T103 = T67[35:32];
  assign T104 = {T108, T105};
  assign T105 = T106;
  assign T106 = T107 != 4'h0;
  assign T107 = T67[39:36];
  assign T108 = T109;
  assign T109 = T110 != 4'h0;
  assign T110 = T67[43:40];
  assign T111 = {T119, T112};
  assign T112 = {T116, T113};
  assign T113 = T114;
  assign T114 = T115 != 4'h0;
  assign T115 = T67[47:44];
  assign T116 = T117;
  assign T117 = T118 != 4'h0;
  assign T118 = T67[51:48];
  assign T119 = T120;
  assign T120 = T121 != 2'h0;
  assign T121 = T67[53:52];
  assign T122 = T123 != 3'h0;
  assign T123 = mainAlignedSigC[2:0];
  assign mainAlignedSigC = $signed(T124) >>> CAlignDist;
  assign T124 = T125;
  assign T125 = {T127, T126};
  assign T126 = 111'h0 - T200;
  assign T200 = {110'h0, doSubMags};
  assign T127 = doSubMags ? T128 : rawC_sig;
  assign T128 = ~ rawC_sig;
  assign T129 = T131 & T130;
  assign T130 = reduced4CExtra ^ 1'h1;
  assign T131 = T132 == 3'h7;
  assign T132 = mainAlignedSigC[2:0];
  assign doSubMags = T134 ^ T133;
  assign T133 = io_op[0];
  assign T134 = signProd ^ rawC_sign;
  assign rawC_sign = T135;
  assign T135 = io_c[64];
  assign signProd = T137 ^ T136;
  assign T136 = io_op[1];
  assign T137 = rawA_sign ^ rawB_sign;
  assign rawB_sign = T138;
  assign T138 = io_b[64];
  assign rawA_sign = T139;
  assign T139 = io_a[64];
  assign T140 = $signed(mainAlignedSigC) >>> 2'h3;
  assign io_toPostMul_highAlignedSigC = T141;
  assign T141 = alignedSigC[161:107];
  assign io_toPostMul_CDom_CAlignDist = T142;
  assign T142 = CAlignDist[5:0];
  assign io_toPostMul_CIsDominant = CIsDominant;
  assign CIsDominant = T145 & T143;
  assign T143 = isMinCAlign | T144;
  assign T144 = posNatCAlignDist <= 13'h35;
  assign T145 = rawC_isZero ^ 1'h1;
  assign rawC_isZero = T72;
  assign io_toPostMul_doSubMags = doSubMags;
  assign io_toPostMul_sExpSum = T201;
  assign T201 = T146[12:0];
  assign T146 = CIsDominant ? T202 : T147;
  assign T147 = sExpAlignedProd - 14'h35;
  assign T202 = {T203, rawC_sExp};
  assign T203 = rawC_sExp[12];
  assign io_toPostMul_isZeroC = rawC_isZero;
  assign io_toPostMul_isInfC = rawC_isInf;
  assign rawC_isInf = T148;
  assign T148 = T151 & T149;
  assign T149 = T150 ^ 1'h1;
  assign T150 = T15[9];
  assign T151 = T152 == 2'h3;
  assign T152 = T15[11:10];
  assign io_toPostMul_isNaNC = rawC_isNaN;
  assign rawC_isNaN = T153;
  assign T153 = T151 & T154;
  assign T154 = T15[9];
  assign io_toPostMul_signProd = signProd;
  assign io_toPostMul_isZeroB = rawB_isZero;
  assign io_toPostMul_isInfB = rawB_isInf;
  assign rawB_isInf = T155;
  assign T155 = T158 & T156;
  assign T156 = T157 ^ 1'h1;
  assign T157 = T19[9];
  assign T158 = T159 == 2'h3;
  assign T159 = T19[11:10];
  assign io_toPostMul_isZeroA = rawA_isZero;
  assign io_toPostMul_isInfA = rawA_isInf;
  assign rawA_isInf = T160;
  assign T160 = T163 & T161;
  assign T161 = T162 ^ 1'h1;
  assign T162 = T22[9];
  assign T163 = T164 == 2'h3;
  assign T164 = T22[11:10];
  assign io_toPostMul_isNaNAOrB = T165;
  assign T165 = rawA_isNaN | rawB_isNaN;
  assign rawB_isNaN = T166;
  assign T166 = T158 & T167;
  assign T167 = T19[9];
  assign rawA_isNaN = T168;
  assign T168 = T163 & T169;
  assign T169 = T22[9];
  assign io_toPostMul_isSigNaNAny = T170;
  assign T170 = T174 | T171;
  assign T171 = rawC_isNaN & T172;
  assign T172 = T173 ^ 1'h1;
  assign T173 = rawC_sig[51];
  assign T174 = T182 | T175;
  assign T175 = rawB_isNaN & T176;
  assign T176 = T177 ^ 1'h1;
  assign T177 = rawB_sig[51];
  assign rawB_sig = T178;
  assign T178 = {1'h0, T179};
  assign T179 = {T181, T180};
  assign T180 = io_b[51:0];
  assign T181 = T26 ^ 1'h1;
  assign T182 = rawA_isNaN & T183;
  assign T183 = T184 ^ 1'h1;
  assign T184 = rawA_sig[51];
  assign rawA_sig = T185;
  assign T185 = {1'h0, T186};
  assign T186 = {T188, T187};
  assign T187 = io_a[51:0];
  assign T188 = T28 ^ 1'h1;
  assign io_mulAddC = T189;
  assign T189 = alignedSigC[106:1];
  assign io_mulAddB = T204;
  assign T204 = rawB_sig[52:0];
  assign io_mulAddA = T205;
  assign T205 = rawA_sig[52:0];
endmodule

module MulAddRecFNToRaw_postMul(
    input  io_fromPreMul_isSigNaNAny,
    input  io_fromPreMul_isNaNAOrB,
    input  io_fromPreMul_isInfA,
    input  io_fromPreMul_isZeroA,
    input  io_fromPreMul_isInfB,
    input  io_fromPreMul_isZeroB,
    input  io_fromPreMul_signProd,
    input  io_fromPreMul_isNaNC,
    input  io_fromPreMul_isInfC,
    input  io_fromPreMul_isZeroC,
    input [12:0] io_fromPreMul_sExpSum,
    input  io_fromPreMul_doSubMags,
    input  io_fromPreMul_CIsDominant,
    input [5:0] io_fromPreMul_CDom_CAlignDist,
    input [54:0] io_fromPreMul_highAlignedSigC,
    input  io_fromPreMul_bit0AlignedSigC,
    input [106:0] io_mulAddResult,
    input [2:0] io_roundingMode,
    output io_invalidExc,
    output io_rawOut_isNaN,
    output io_rawOut_isInf,
    output io_rawOut_isZero,
    output io_rawOut_sign,
    output[12:0] io_rawOut_sExp,
    output[55:0] io_rawOut_sig
);

  wire[55:0] T0;
  wire[55:0] notCDom_sig;
  wire T1;
  wire notCDom_reduced4SigExtra;
  wire[13:0] T2;
  wire[13:0] T561;
  wire[12:0] T3;
  wire[4:0] T4;
  wire T5;
  wire[4:0] T6;
  wire[12:0] T7;
  wire[32:0] T8;
  wire[4:0] T9;
  wire[4:0] T10;
  wire[5:0] T562;
  wire[5:0] T563;
  wire[5:0] T564;
  wire[5:0] T565;
  wire[5:0] T566;
  wire[5:0] T567;
  wire[5:0] T568;
  wire[5:0] T569;
  wire[5:0] T570;
  wire[5:0] T571;
  wire[5:0] T572;
  wire[5:0] T573;
  wire[5:0] T574;
  wire[5:0] T575;
  wire[5:0] T576;
  wire[5:0] T577;
  wire[5:0] T578;
  wire[5:0] T579;
  wire[5:0] T580;
  wire[5:0] T581;
  wire[5:0] T582;
  wire[5:0] T583;
  wire[5:0] T584;
  wire[5:0] T585;
  wire[5:0] T586;
  wire[5:0] T587;
  wire[5:0] T588;
  wire[5:0] T589;
  wire[5:0] T590;
  wire[5:0] T591;
  wire[5:0] T592;
  wire[5:0] T593;
  wire[5:0] T594;
  wire[5:0] T595;
  wire[5:0] T596;
  wire[5:0] T597;
  wire[5:0] T598;
  wire[5:0] T599;
  wire[5:0] T600;
  wire[5:0] T601;
  wire[5:0] T602;
  wire[5:0] T603;
  wire[5:0] T604;
  wire[5:0] T605;
  wire[5:0] T606;
  wire[5:0] T607;
  wire[5:0] T608;
  wire[5:0] T609;
  wire[5:0] T610;
  wire[5:0] T611;
  wire[5:0] T612;
  wire[5:0] T613;
  wire[5:0] T614;
  wire[5:0] T615;
  wire T616;
  wire[54:0] T11;
  wire[22:0] T12;
  wire[6:0] T13;
  wire[2:0] T14;
  wire T15;
  wire[2:0] T16;
  wire[6:0] T17;
  wire[22:0] T18;
  wire[54:0] notCDom_reduced2AbsSigSum;
  wire[54:0] T19;
  wire[27:0] T20;
  wire[13:0] T21;
  wire[6:0] T22;
  wire[3:0] T23;
  wire[1:0] T24;
  wire T25;
  wire T26;
  wire[1:0] T27;
  wire[108:0] notCDom_absSigSum;
  wire[108:0] T28;
  wire[108:0] T617;
  wire[108:0] T29;
  wire[161:0] sigSum;
  wire[106:0] T30;
  wire[105:0] T31;
  wire[54:0] T32;
  wire[54:0] T33;
  wire T34;
  wire[108:0] T35;
  wire[108:0] T36;
  wire notCDom_signSigSum;
  wire T37;
  wire T38;
  wire[1:0] T39;
  wire[1:0] T40;
  wire T41;
  wire T42;
  wire[1:0] T43;
  wire T44;
  wire T45;
  wire[1:0] T46;
  wire[2:0] T47;
  wire[1:0] T48;
  wire T49;
  wire T50;
  wire[1:0] T51;
  wire T52;
  wire T53;
  wire[1:0] T54;
  wire T55;
  wire T56;
  wire[1:0] T57;
  wire[6:0] T58;
  wire[3:0] T59;
  wire[1:0] T60;
  wire T61;
  wire T62;
  wire[1:0] T63;
  wire T64;
  wire T65;
  wire[1:0] T66;
  wire[1:0] T67;
  wire T68;
  wire T69;
  wire[1:0] T70;
  wire T71;
  wire T72;
  wire[1:0] T73;
  wire[2:0] T74;
  wire[1:0] T75;
  wire T76;
  wire T77;
  wire[1:0] T78;
  wire T79;
  wire T80;
  wire[1:0] T81;
  wire T82;
  wire T83;
  wire[1:0] T84;
  wire[13:0] T85;
  wire[6:0] T86;
  wire[3:0] T87;
  wire[1:0] T88;
  wire T89;
  wire T90;
  wire[1:0] T91;
  wire T92;
  wire T93;
  wire[1:0] T94;
  wire[1:0] T95;
  wire T96;
  wire T97;
  wire[1:0] T98;
  wire T99;
  wire T100;
  wire[1:0] T101;
  wire[2:0] T102;
  wire[1:0] T103;
  wire T104;
  wire T105;
  wire[1:0] T106;
  wire T107;
  wire T108;
  wire[1:0] T109;
  wire T110;
  wire T111;
  wire[1:0] T112;
  wire[6:0] T113;
  wire[3:0] T114;
  wire[1:0] T115;
  wire T116;
  wire T117;
  wire[1:0] T118;
  wire T119;
  wire T120;
  wire[1:0] T121;
  wire[1:0] T122;
  wire T123;
  wire T124;
  wire[1:0] T125;
  wire T126;
  wire T127;
  wire[1:0] T128;
  wire[2:0] T129;
  wire[1:0] T130;
  wire T131;
  wire T132;
  wire[1:0] T133;
  wire T134;
  wire T135;
  wire[1:0] T136;
  wire T137;
  wire T138;
  wire[1:0] T139;
  wire[26:0] T140;
  wire[13:0] T141;
  wire[6:0] T142;
  wire[3:0] T143;
  wire[1:0] T144;
  wire T145;
  wire T146;
  wire[1:0] T147;
  wire T148;
  wire T149;
  wire[1:0] T150;
  wire[1:0] T151;
  wire T152;
  wire T153;
  wire[1:0] T154;
  wire T155;
  wire T156;
  wire[1:0] T157;
  wire[2:0] T158;
  wire[1:0] T159;
  wire T160;
  wire T161;
  wire[1:0] T162;
  wire T163;
  wire T164;
  wire[1:0] T165;
  wire T166;
  wire T167;
  wire[1:0] T168;
  wire[6:0] T169;
  wire[3:0] T170;
  wire[1:0] T171;
  wire T172;
  wire T173;
  wire[1:0] T174;
  wire T175;
  wire T176;
  wire[1:0] T177;
  wire[1:0] T178;
  wire T179;
  wire T180;
  wire[1:0] T181;
  wire T182;
  wire T183;
  wire[1:0] T184;
  wire[2:0] T185;
  wire[1:0] T186;
  wire T187;
  wire T188;
  wire[1:0] T189;
  wire T190;
  wire T191;
  wire[1:0] T192;
  wire T193;
  wire T194;
  wire[1:0] T195;
  wire[12:0] T196;
  wire[6:0] T197;
  wire[3:0] T198;
  wire[1:0] T199;
  wire T200;
  wire T201;
  wire[1:0] T202;
  wire T203;
  wire T204;
  wire[1:0] T205;
  wire[1:0] T206;
  wire T207;
  wire T208;
  wire[1:0] T209;
  wire T210;
  wire T211;
  wire[1:0] T212;
  wire[2:0] T213;
  wire[1:0] T214;
  wire T215;
  wire T216;
  wire[1:0] T217;
  wire T218;
  wire T219;
  wire[1:0] T220;
  wire T221;
  wire T222;
  wire[1:0] T223;
  wire[5:0] T224;
  wire[2:0] T225;
  wire[1:0] T226;
  wire T227;
  wire T228;
  wire[1:0] T229;
  wire T230;
  wire T231;
  wire[1:0] T232;
  wire T233;
  wire T234;
  wire[1:0] T235;
  wire[2:0] T236;
  wire[1:0] T237;
  wire T238;
  wire T239;
  wire[1:0] T240;
  wire T241;
  wire T242;
  wire[1:0] T243;
  wire T244;
  wire T245;
  wire T246;
  wire[1:0] T247;
  wire T248;
  wire[1:0] T249;
  wire T250;
  wire[3:0] T251;
  wire[1:0] T252;
  wire T253;
  wire[1:0] T254;
  wire[3:0] T255;
  wire T256;
  wire[1:0] T257;
  wire T258;
  wire[1:0] T259;
  wire T260;
  wire[15:0] T261;
  wire[15:0] T262;
  wire[15:0] T263;
  wire[14:0] T264;
  wire[15:0] T265;
  wire[15:0] T266;
  wire[15:0] T267;
  wire[13:0] T268;
  wire[15:0] T269;
  wire[15:0] T270;
  wire[15:0] T271;
  wire[11:0] T272;
  wire[15:0] T273;
  wire[15:0] T274;
  wire[15:0] T275;
  wire[7:0] T276;
  wire[15:0] T277;
  wire[15:0] T278;
  wire[15:0] T618;
  wire[7:0] T279;
  wire[15:0] T280;
  wire[15:0] T619;
  wire[11:0] T281;
  wire[15:0] T282;
  wire[15:0] T620;
  wire[13:0] T283;
  wire[15:0] T284;
  wire[15:0] T621;
  wire[14:0] T285;
  wire[31:0] T286;
  wire[31:0] T287;
  wire[31:0] T288;
  wire[30:0] T289;
  wire[31:0] T290;
  wire[31:0] T291;
  wire[31:0] T292;
  wire[29:0] T293;
  wire[31:0] T294;
  wire[31:0] T295;
  wire[31:0] T296;
  wire[27:0] T297;
  wire[31:0] T298;
  wire[31:0] T299;
  wire[31:0] T300;
  wire[23:0] T301;
  wire[31:0] T302;
  wire[31:0] T303;
  wire[31:0] T304;
  wire[15:0] T305;
  wire[31:0] T306;
  wire[31:0] T307;
  wire[31:0] T622;
  wire[15:0] T308;
  wire[31:0] T309;
  wire[31:0] T623;
  wire[23:0] T310;
  wire[31:0] T311;
  wire[31:0] T624;
  wire[27:0] T312;
  wire[31:0] T313;
  wire[31:0] T625;
  wire[29:0] T314;
  wire[31:0] T315;
  wire[31:0] T626;
  wire[30:0] T316;
  wire T627;
  wire T628;
  wire T629;
  wire T630;
  wire T631;
  wire T632;
  wire T633;
  wire T634;
  wire T635;
  wire T636;
  wire T637;
  wire T638;
  wire T639;
  wire T640;
  wire T641;
  wire T642;
  wire T643;
  wire T644;
  wire T645;
  wire T646;
  wire T647;
  wire T648;
  wire T649;
  wire T650;
  wire T651;
  wire T652;
  wire T653;
  wire T654;
  wire T655;
  wire T656;
  wire T657;
  wire T658;
  wire T659;
  wire T660;
  wire T661;
  wire T662;
  wire T663;
  wire T664;
  wire T665;
  wire T666;
  wire T667;
  wire T668;
  wire T669;
  wire T670;
  wire T671;
  wire T672;
  wire T673;
  wire T674;
  wire T675;
  wire T676;
  wire T677;
  wire T678;
  wire T679;
  wire[3:0] T317;
  wire[1:0] T318;
  wire T319;
  wire[1:0] T320;
  wire[3:0] T321;
  wire T322;
  wire[1:0] T323;
  wire T324;
  wire[1:0] T325;
  wire T326;
  wire[7:0] T327;
  wire[7:0] T328;
  wire[7:0] T329;
  wire[6:0] T330;
  wire[7:0] T331;
  wire[7:0] T332;
  wire[7:0] T333;
  wire[5:0] T334;
  wire[7:0] T335;
  wire[7:0] T336;
  wire[7:0] T337;
  wire[3:0] T338;
  wire[7:0] T339;
  wire[7:0] T340;
  wire[7:0] T680;
  wire[3:0] T341;
  wire[7:0] T342;
  wire[7:0] T681;
  wire[5:0] T343;
  wire[7:0] T344;
  wire[7:0] T682;
  wire[6:0] T345;
  wire[13:0] T346;
  wire[13:0] T347;
  wire[6:0] T348;
  wire[3:0] T349;
  wire[1:0] T350;
  wire T351;
  wire T352;
  wire[1:0] T353;
  wire[26:0] T354;
  wire[26:0] T355;
  wire T356;
  wire T357;
  wire[1:0] T358;
  wire[1:0] T359;
  wire T360;
  wire T361;
  wire[1:0] T362;
  wire T363;
  wire T364;
  wire[1:0] T365;
  wire[2:0] T366;
  wire[1:0] T367;
  wire T368;
  wire T369;
  wire[1:0] T370;
  wire T371;
  wire T372;
  wire[1:0] T373;
  wire T374;
  wire T375;
  wire[1:0] T376;
  wire[6:0] T377;
  wire[3:0] T378;
  wire[1:0] T379;
  wire T380;
  wire T381;
  wire[1:0] T382;
  wire T383;
  wire T384;
  wire[1:0] T385;
  wire[1:0] T386;
  wire T387;
  wire T388;
  wire[1:0] T389;
  wire T390;
  wire T391;
  wire[1:0] T392;
  wire[2:0] T393;
  wire[1:0] T394;
  wire T395;
  wire T396;
  wire[1:0] T397;
  wire T398;
  wire T399;
  wire[1:0] T400;
  wire T401;
  wire T402;
  wire T403;
  wire T404;
  wire[2:0] T405;
  wire[57:0] notCDom_mainSig;
  wire[235:0] T406;
  wire[6:0] notCDom_nearNormDist;
  wire[54:0] T407;
  wire[55:0] CDom_sig;
  wire T408;
  wire CDom_absSigSumExtra;
  wire T409;
  wire[53:0] T410;
  wire T411;
  wire[52:0] T412;
  wire[52:0] T413;
  wire T414;
  wire CDom_reduced4SigExtra;
  wire[13:0] T415;
  wire[13:0] T683;
  wire[12:0] T416;
  wire[4:0] T417;
  wire T418;
  wire[4:0] T419;
  wire[12:0] T420;
  wire[16:0] T421;
  wire[3:0] T422;
  wire[3:0] T423;
  wire[3:0] T424;
  wire[1:0] T425;
  wire T426;
  wire[1:0] T427;
  wire[3:0] T428;
  wire T429;
  wire[1:0] T430;
  wire T431;
  wire[1:0] T432;
  wire T433;
  wire[7:0] T434;
  wire[7:0] T435;
  wire[7:0] T436;
  wire[6:0] T437;
  wire[7:0] T438;
  wire[7:0] T439;
  wire[7:0] T440;
  wire[5:0] T441;
  wire[7:0] T442;
  wire[7:0] T443;
  wire[7:0] T444;
  wire[3:0] T445;
  wire[7:0] T446;
  wire[7:0] T447;
  wire[7:0] T684;
  wire[3:0] T448;
  wire[7:0] T449;
  wire[7:0] T685;
  wire[5:0] T450;
  wire[7:0] T451;
  wire[7:0] T686;
  wire[6:0] T452;
  wire[13:0] T453;
  wire[13:0] T454;
  wire[6:0] T455;
  wire[3:0] T456;
  wire[1:0] T457;
  wire T458;
  wire T459;
  wire[3:0] T460;
  wire[54:0] T461;
  wire[52:0] T462;
  wire[107:0] CDom_absSigSum;
  wire[107:0] T463;
  wire[106:0] T464;
  wire[104:0] T465;
  wire[1:0] T466;
  wire[107:0] T467;
  wire[107:0] T468;
  wire T469;
  wire T470;
  wire[3:0] T471;
  wire[1:0] T472;
  wire T473;
  wire T474;
  wire[3:0] T475;
  wire T476;
  wire T477;
  wire[3:0] T478;
  wire[2:0] T479;
  wire[1:0] T480;
  wire T481;
  wire T482;
  wire[3:0] T483;
  wire T484;
  wire T485;
  wire[3:0] T486;
  wire T487;
  wire T488;
  wire[3:0] T489;
  wire[6:0] T490;
  wire[3:0] T491;
  wire[1:0] T492;
  wire T493;
  wire T494;
  wire[3:0] T495;
  wire T496;
  wire T497;
  wire[3:0] T498;
  wire[1:0] T499;
  wire T500;
  wire T501;
  wire[3:0] T502;
  wire T503;
  wire T504;
  wire[3:0] T505;
  wire[2:0] T506;
  wire[1:0] T507;
  wire T508;
  wire T509;
  wire[3:0] T510;
  wire T511;
  wire T512;
  wire[3:0] T513;
  wire T514;
  wire T515;
  wire[2:0] T516;
  wire T517;
  wire[2:0] T518;
  wire[57:0] CDom_mainSig;
  wire[170:0] T519;
  wire[54:0] T520;
  wire[12:0] T521;
  wire[12:0] notCDom_sExp;
  wire[12:0] T687;
  wire[7:0] T522;
  wire[7:0] T523;
  wire[4:0] T688;
  wire T689;
  wire[12:0] CDom_sExp;
  wire[12:0] T690;
  wire[1:0] T524;
  wire[1:0] T525;
  wire[10:0] T691;
  wire T692;
  wire T526;
  wire T527;
  wire T528;
  wire notCDom_sign;
  wire T529;
  wire roundingMode_min;
  wire notCDom_completeCancellation;
  wire[1:0] T530;
  wire CDom_sign;
  wire T531;
  wire T532;
  wire notNaN_addZeros;
  wire T533;
  wire T534;
  wire notNaN_isInfOut;
  wire notNaN_isInfProd;
  wire T535;
  wire T536;
  wire T537;
  wire T538;
  wire T539;
  wire T540;
  wire T541;
  wire T542;
  wire T543;
  wire T544;
  wire T545;
  wire T546;
  wire T547;
  wire T548;
  wire T549;
  wire T550;
  wire T551;
  wire T552;
  wire T553;
  wire T554;
  wire T555;
  wire T556;
  wire T557;
  wire T558;
  wire T559;
  wire T560;


  assign io_rawOut_sig = T0;
  assign T0 = io_fromPreMul_CIsDominant ? CDom_sig : notCDom_sig;
  assign notCDom_sig = {T407, T1};
  assign T1 = T404 | notCDom_reduced4SigExtra;
  assign notCDom_reduced4SigExtra = T2 != 14'h0;
  assign T2 = T346 & T561;
  assign T561 = {1'h0, T3};
  assign T3 = {T327, T4};
  assign T4 = {T317, T5};
  assign T5 = T6[4];
  assign T6 = T7[12:8];
  assign T7 = T8[13:1];
  assign T8 = $signed(33'h100000000) >>> T9;
  assign T9 = ~ T10;
  assign T10 = T562 >> 1'h1;
  assign T562 = T679 ? 1'h0 : T563;
  assign T563 = T678 ? 1'h1 : T564;
  assign T564 = T677 ? 2'h2 : T565;
  assign T565 = T676 ? 2'h3 : T566;
  assign T566 = T675 ? 3'h4 : T567;
  assign T567 = T674 ? 3'h5 : T568;
  assign T568 = T673 ? 3'h6 : T569;
  assign T569 = T672 ? 3'h7 : T570;
  assign T570 = T671 ? 4'h8 : T571;
  assign T571 = T670 ? 4'h9 : T572;
  assign T572 = T669 ? 4'ha : T573;
  assign T573 = T668 ? 4'hb : T574;
  assign T574 = T667 ? 4'hc : T575;
  assign T575 = T666 ? 4'hd : T576;
  assign T576 = T665 ? 4'he : T577;
  assign T577 = T664 ? 4'hf : T578;
  assign T578 = T663 ? 5'h10 : T579;
  assign T579 = T662 ? 5'h11 : T580;
  assign T580 = T661 ? 5'h12 : T581;
  assign T581 = T660 ? 5'h13 : T582;
  assign T582 = T659 ? 5'h14 : T583;
  assign T583 = T658 ? 5'h15 : T584;
  assign T584 = T657 ? 5'h16 : T585;
  assign T585 = T656 ? 5'h17 : T586;
  assign T586 = T655 ? 5'h18 : T587;
  assign T587 = T654 ? 5'h19 : T588;
  assign T588 = T653 ? 5'h1a : T589;
  assign T589 = T652 ? 5'h1b : T590;
  assign T590 = T651 ? 5'h1c : T591;
  assign T591 = T650 ? 5'h1d : T592;
  assign T592 = T649 ? 5'h1e : T593;
  assign T593 = T648 ? 5'h1f : T594;
  assign T594 = T647 ? 6'h20 : T595;
  assign T595 = T646 ? 6'h21 : T596;
  assign T596 = T645 ? 6'h22 : T597;
  assign T597 = T644 ? 6'h23 : T598;
  assign T598 = T643 ? 6'h24 : T599;
  assign T599 = T642 ? 6'h25 : T600;
  assign T600 = T641 ? 6'h26 : T601;
  assign T601 = T640 ? 6'h27 : T602;
  assign T602 = T639 ? 6'h28 : T603;
  assign T603 = T638 ? 6'h29 : T604;
  assign T604 = T637 ? 6'h2a : T605;
  assign T605 = T636 ? 6'h2b : T606;
  assign T606 = T635 ? 6'h2c : T607;
  assign T607 = T634 ? 6'h2d : T608;
  assign T608 = T633 ? 6'h2e : T609;
  assign T609 = T632 ? 6'h2f : T610;
  assign T610 = T631 ? 6'h30 : T611;
  assign T611 = T630 ? 6'h31 : T612;
  assign T612 = T629 ? 6'h32 : T613;
  assign T613 = T628 ? 6'h33 : T614;
  assign T614 = T627 ? 6'h34 : T615;
  assign T615 = T616 ? 6'h35 : 6'h36;
  assign T616 = T11[53];
  assign T11 = {T286, T12};
  assign T12 = {T261, T13};
  assign T13 = {T251, T14};
  assign T14 = {T247, T15};
  assign T15 = T16[2];
  assign T16 = T17[6:4];
  assign T17 = T18[22:16];
  assign T18 = notCDom_reduced2AbsSigSum[54:32];
  assign notCDom_reduced2AbsSigSum = T19;
  assign T19 = {T140, T20};
  assign T20 = {T85, T21};
  assign T21 = {T58, T22};
  assign T22 = {T47, T23};
  assign T23 = {T40, T24};
  assign T24 = {T37, T25};
  assign T25 = T26;
  assign T26 = T27 != 2'h0;
  assign T27 = notCDom_absSigSum[1:0];
  assign notCDom_absSigSum = notCDom_signSigSum ? T35 : T28;
  assign T28 = T29 + T617;
  assign T617 = {108'h0, io_fromPreMul_doSubMags};
  assign T29 = sigSum[108:0];
  assign sigSum = {T32, T30};
  assign T30 = {T31, io_fromPreMul_bit0AlignedSigC};
  assign T31 = io_mulAddResult[105:0];
  assign T32 = T34 ? T33 : io_fromPreMul_highAlignedSigC;
  assign T33 = io_fromPreMul_highAlignedSigC + 55'h1;
  assign T34 = io_mulAddResult[106];
  assign T35 = ~ T36;
  assign T36 = sigSum[108:0];
  assign notCDom_signSigSum = sigSum[109];
  assign T37 = T38;
  assign T38 = T39 != 2'h0;
  assign T39 = notCDom_absSigSum[3:2];
  assign T40 = {T44, T41};
  assign T41 = T42;
  assign T42 = T43 != 2'h0;
  assign T43 = notCDom_absSigSum[5:4];
  assign T44 = T45;
  assign T45 = T46 != 2'h0;
  assign T46 = notCDom_absSigSum[7:6];
  assign T47 = {T55, T48};
  assign T48 = {T52, T49};
  assign T49 = T50;
  assign T50 = T51 != 2'h0;
  assign T51 = notCDom_absSigSum[9:8];
  assign T52 = T53;
  assign T53 = T54 != 2'h0;
  assign T54 = notCDom_absSigSum[11:10];
  assign T55 = T56;
  assign T56 = T57 != 2'h0;
  assign T57 = notCDom_absSigSum[13:12];
  assign T58 = {T74, T59};
  assign T59 = {T67, T60};
  assign T60 = {T64, T61};
  assign T61 = T62;
  assign T62 = T63 != 2'h0;
  assign T63 = notCDom_absSigSum[15:14];
  assign T64 = T65;
  assign T65 = T66 != 2'h0;
  assign T66 = notCDom_absSigSum[17:16];
  assign T67 = {T71, T68};
  assign T68 = T69;
  assign T69 = T70 != 2'h0;
  assign T70 = notCDom_absSigSum[19:18];
  assign T71 = T72;
  assign T72 = T73 != 2'h0;
  assign T73 = notCDom_absSigSum[21:20];
  assign T74 = {T82, T75};
  assign T75 = {T79, T76};
  assign T76 = T77;
  assign T77 = T78 != 2'h0;
  assign T78 = notCDom_absSigSum[23:22];
  assign T79 = T80;
  assign T80 = T81 != 2'h0;
  assign T81 = notCDom_absSigSum[25:24];
  assign T82 = T83;
  assign T83 = T84 != 2'h0;
  assign T84 = notCDom_absSigSum[27:26];
  assign T85 = {T113, T86};
  assign T86 = {T102, T87};
  assign T87 = {T95, T88};
  assign T88 = {T92, T89};
  assign T89 = T90;
  assign T90 = T91 != 2'h0;
  assign T91 = notCDom_absSigSum[29:28];
  assign T92 = T93;
  assign T93 = T94 != 2'h0;
  assign T94 = notCDom_absSigSum[31:30];
  assign T95 = {T99, T96};
  assign T96 = T97;
  assign T97 = T98 != 2'h0;
  assign T98 = notCDom_absSigSum[33:32];
  assign T99 = T100;
  assign T100 = T101 != 2'h0;
  assign T101 = notCDom_absSigSum[35:34];
  assign T102 = {T110, T103};
  assign T103 = {T107, T104};
  assign T104 = T105;
  assign T105 = T106 != 2'h0;
  assign T106 = notCDom_absSigSum[37:36];
  assign T107 = T108;
  assign T108 = T109 != 2'h0;
  assign T109 = notCDom_absSigSum[39:38];
  assign T110 = T111;
  assign T111 = T112 != 2'h0;
  assign T112 = notCDom_absSigSum[41:40];
  assign T113 = {T129, T114};
  assign T114 = {T122, T115};
  assign T115 = {T119, T116};
  assign T116 = T117;
  assign T117 = T118 != 2'h0;
  assign T118 = notCDom_absSigSum[43:42];
  assign T119 = T120;
  assign T120 = T121 != 2'h0;
  assign T121 = notCDom_absSigSum[45:44];
  assign T122 = {T126, T123};
  assign T123 = T124;
  assign T124 = T125 != 2'h0;
  assign T125 = notCDom_absSigSum[47:46];
  assign T126 = T127;
  assign T127 = T128 != 2'h0;
  assign T128 = notCDom_absSigSum[49:48];
  assign T129 = {T137, T130};
  assign T130 = {T134, T131};
  assign T131 = T132;
  assign T132 = T133 != 2'h0;
  assign T133 = notCDom_absSigSum[51:50];
  assign T134 = T135;
  assign T135 = T136 != 2'h0;
  assign T136 = notCDom_absSigSum[53:52];
  assign T137 = T138;
  assign T138 = T139 != 2'h0;
  assign T139 = notCDom_absSigSum[55:54];
  assign T140 = {T196, T141};
  assign T141 = {T169, T142};
  assign T142 = {T158, T143};
  assign T143 = {T151, T144};
  assign T144 = {T148, T145};
  assign T145 = T146;
  assign T146 = T147 != 2'h0;
  assign T147 = notCDom_absSigSum[57:56];
  assign T148 = T149;
  assign T149 = T150 != 2'h0;
  assign T150 = notCDom_absSigSum[59:58];
  assign T151 = {T155, T152};
  assign T152 = T153;
  assign T153 = T154 != 2'h0;
  assign T154 = notCDom_absSigSum[61:60];
  assign T155 = T156;
  assign T156 = T157 != 2'h0;
  assign T157 = notCDom_absSigSum[63:62];
  assign T158 = {T166, T159};
  assign T159 = {T163, T160};
  assign T160 = T161;
  assign T161 = T162 != 2'h0;
  assign T162 = notCDom_absSigSum[65:64];
  assign T163 = T164;
  assign T164 = T165 != 2'h0;
  assign T165 = notCDom_absSigSum[67:66];
  assign T166 = T167;
  assign T167 = T168 != 2'h0;
  assign T168 = notCDom_absSigSum[69:68];
  assign T169 = {T185, T170};
  assign T170 = {T178, T171};
  assign T171 = {T175, T172};
  assign T172 = T173;
  assign T173 = T174 != 2'h0;
  assign T174 = notCDom_absSigSum[71:70];
  assign T175 = T176;
  assign T176 = T177 != 2'h0;
  assign T177 = notCDom_absSigSum[73:72];
  assign T178 = {T182, T179};
  assign T179 = T180;
  assign T180 = T181 != 2'h0;
  assign T181 = notCDom_absSigSum[75:74];
  assign T182 = T183;
  assign T183 = T184 != 2'h0;
  assign T184 = notCDom_absSigSum[77:76];
  assign T185 = {T193, T186};
  assign T186 = {T190, T187};
  assign T187 = T188;
  assign T188 = T189 != 2'h0;
  assign T189 = notCDom_absSigSum[79:78];
  assign T190 = T191;
  assign T191 = T192 != 2'h0;
  assign T192 = notCDom_absSigSum[81:80];
  assign T193 = T194;
  assign T194 = T195 != 2'h0;
  assign T195 = notCDom_absSigSum[83:82];
  assign T196 = {T224, T197};
  assign T197 = {T213, T198};
  assign T198 = {T206, T199};
  assign T199 = {T203, T200};
  assign T200 = T201;
  assign T201 = T202 != 2'h0;
  assign T202 = notCDom_absSigSum[85:84];
  assign T203 = T204;
  assign T204 = T205 != 2'h0;
  assign T205 = notCDom_absSigSum[87:86];
  assign T206 = {T210, T207};
  assign T207 = T208;
  assign T208 = T209 != 2'h0;
  assign T209 = notCDom_absSigSum[89:88];
  assign T210 = T211;
  assign T211 = T212 != 2'h0;
  assign T212 = notCDom_absSigSum[91:90];
  assign T213 = {T221, T214};
  assign T214 = {T218, T215};
  assign T215 = T216;
  assign T216 = T217 != 2'h0;
  assign T217 = notCDom_absSigSum[93:92];
  assign T218 = T219;
  assign T219 = T220 != 2'h0;
  assign T220 = notCDom_absSigSum[95:94];
  assign T221 = T222;
  assign T222 = T223 != 2'h0;
  assign T223 = notCDom_absSigSum[97:96];
  assign T224 = {T236, T225};
  assign T225 = {T233, T226};
  assign T226 = {T230, T227};
  assign T227 = T228;
  assign T228 = T229 != 2'h0;
  assign T229 = notCDom_absSigSum[99:98];
  assign T230 = T231;
  assign T231 = T232 != 2'h0;
  assign T232 = notCDom_absSigSum[101:100];
  assign T233 = T234;
  assign T234 = T235 != 2'h0;
  assign T235 = notCDom_absSigSum[103:102];
  assign T236 = {T244, T237};
  assign T237 = {T241, T238};
  assign T238 = T239;
  assign T239 = T240 != 2'h0;
  assign T240 = notCDom_absSigSum[105:104];
  assign T241 = T242;
  assign T242 = T243 != 2'h0;
  assign T243 = notCDom_absSigSum[107:106];
  assign T244 = T245;
  assign T245 = T246 != 1'h0;
  assign T246 = notCDom_absSigSum[108];
  assign T247 = {T250, T248};
  assign T248 = T249[1];
  assign T249 = T16[1:0];
  assign T250 = T249[0];
  assign T251 = {T257, T252};
  assign T252 = {T256, T253};
  assign T253 = T254[1];
  assign T254 = T255[3:2];
  assign T255 = T17[3:0];
  assign T256 = T254[0];
  assign T257 = {T260, T258};
  assign T258 = T259[1];
  assign T259 = T255[1:0];
  assign T260 = T259[0];
  assign T261 = T284 | T262;
  assign T262 = T263 & 16'haaaa;
  assign T263 = T264 << 1'h1;
  assign T264 = T265[14:0];
  assign T265 = T282 | T266;
  assign T266 = T267 & 16'hcccc;
  assign T267 = T268 << 2'h2;
  assign T268 = T269[13:0];
  assign T269 = T280 | T270;
  assign T270 = T271 & 16'hf0f0;
  assign T271 = T272 << 3'h4;
  assign T272 = T273[11:0];
  assign T273 = T278 | T274;
  assign T274 = T275 & 16'hff00;
  assign T275 = T276 << 4'h8;
  assign T276 = T277[7:0];
  assign T277 = T18[15:0];
  assign T278 = T618 & 16'hff;
  assign T618 = {8'h0, T279};
  assign T279 = T277 >> 4'h8;
  assign T280 = T619 & 16'hf0f;
  assign T619 = {4'h0, T281};
  assign T281 = T273 >> 3'h4;
  assign T282 = T620 & 16'h3333;
  assign T620 = {2'h0, T283};
  assign T283 = T269 >> 2'h2;
  assign T284 = T621 & 16'h5555;
  assign T621 = {1'h0, T285};
  assign T285 = T265 >> 1'h1;
  assign T286 = T315 | T287;
  assign T287 = T288 & 32'haaaaaaaa;
  assign T288 = T289 << 1'h1;
  assign T289 = T290[30:0];
  assign T290 = T313 | T291;
  assign T291 = T292 & 32'hcccccccc;
  assign T292 = T293 << 2'h2;
  assign T293 = T294[29:0];
  assign T294 = T311 | T295;
  assign T295 = T296 & 32'hf0f0f0f0;
  assign T296 = T297 << 3'h4;
  assign T297 = T298[27:0];
  assign T298 = T309 | T299;
  assign T299 = T300 & 32'hff00ff00;
  assign T300 = T301 << 4'h8;
  assign T301 = T302[23:0];
  assign T302 = T307 | T303;
  assign T303 = T304 & 32'hffff0000;
  assign T304 = T305 << 5'h10;
  assign T305 = T306[15:0];
  assign T306 = notCDom_reduced2AbsSigSum[31:0];
  assign T307 = T622 & 32'hffff;
  assign T622 = {16'h0, T308};
  assign T308 = T306 >> 5'h10;
  assign T309 = T623 & 32'hff00ff;
  assign T623 = {8'h0, T310};
  assign T310 = T302 >> 4'h8;
  assign T311 = T624 & 32'hf0f0f0f;
  assign T624 = {4'h0, T312};
  assign T312 = T298 >> 3'h4;
  assign T313 = T625 & 32'h33333333;
  assign T625 = {2'h0, T314};
  assign T314 = T294 >> 2'h2;
  assign T315 = T626 & 32'h55555555;
  assign T626 = {1'h0, T316};
  assign T316 = T290 >> 1'h1;
  assign T627 = T11[52];
  assign T628 = T11[51];
  assign T629 = T11[50];
  assign T630 = T11[49];
  assign T631 = T11[48];
  assign T632 = T11[47];
  assign T633 = T11[46];
  assign T634 = T11[45];
  assign T635 = T11[44];
  assign T636 = T11[43];
  assign T637 = T11[42];
  assign T638 = T11[41];
  assign T639 = T11[40];
  assign T640 = T11[39];
  assign T641 = T11[38];
  assign T642 = T11[37];
  assign T643 = T11[36];
  assign T644 = T11[35];
  assign T645 = T11[34];
  assign T646 = T11[33];
  assign T647 = T11[32];
  assign T648 = T11[31];
  assign T649 = T11[30];
  assign T650 = T11[29];
  assign T651 = T11[28];
  assign T652 = T11[27];
  assign T653 = T11[26];
  assign T654 = T11[25];
  assign T655 = T11[24];
  assign T656 = T11[23];
  assign T657 = T11[22];
  assign T658 = T11[21];
  assign T659 = T11[20];
  assign T660 = T11[19];
  assign T661 = T11[18];
  assign T662 = T11[17];
  assign T663 = T11[16];
  assign T664 = T11[15];
  assign T665 = T11[14];
  assign T666 = T11[13];
  assign T667 = T11[12];
  assign T668 = T11[11];
  assign T669 = T11[10];
  assign T670 = T11[9];
  assign T671 = T11[8];
  assign T672 = T11[7];
  assign T673 = T11[6];
  assign T674 = T11[5];
  assign T675 = T11[4];
  assign T676 = T11[3];
  assign T677 = T11[2];
  assign T678 = T11[1];
  assign T679 = T11[0];
  assign T317 = {T323, T318};
  assign T318 = {T322, T319};
  assign T319 = T320[1];
  assign T320 = T321[3:2];
  assign T321 = T6[3:0];
  assign T322 = T320[0];
  assign T323 = {T326, T324};
  assign T324 = T325[1];
  assign T325 = T321[1:0];
  assign T326 = T325[0];
  assign T327 = T344 | T328;
  assign T328 = T329 & 8'haa;
  assign T329 = T330 << 1'h1;
  assign T330 = T331[6:0];
  assign T331 = T342 | T332;
  assign T332 = T333 & 8'hcc;
  assign T333 = T334 << 2'h2;
  assign T334 = T335[5:0];
  assign T335 = T340 | T336;
  assign T336 = T337 & 8'hf0;
  assign T337 = T338 << 3'h4;
  assign T338 = T339[3:0];
  assign T339 = T7[7:0];
  assign T340 = T680 & 8'hf;
  assign T680 = {4'h0, T341};
  assign T341 = T339 >> 3'h4;
  assign T342 = T681 & 8'h33;
  assign T681 = {2'h0, T343};
  assign T343 = T335 >> 2'h2;
  assign T344 = T682 & 8'h55;
  assign T682 = {1'h0, T345};
  assign T345 = T331 >> 1'h1;
  assign T346 = T347;
  assign T347 = {T377, T348};
  assign T348 = {T366, T349};
  assign T349 = {T359, T350};
  assign T350 = {T356, T351};
  assign T351 = T352;
  assign T352 = T353 != 2'h0;
  assign T353 = T354[1:0];
  assign T354 = T355 << 1'h0;
  assign T355 = notCDom_reduced2AbsSigSum[26:0];
  assign T356 = T357;
  assign T357 = T358 != 2'h0;
  assign T358 = T354[3:2];
  assign T359 = {T363, T360};
  assign T360 = T361;
  assign T361 = T362 != 2'h0;
  assign T362 = T354[5:4];
  assign T363 = T364;
  assign T364 = T365 != 2'h0;
  assign T365 = T354[7:6];
  assign T366 = {T374, T367};
  assign T367 = {T371, T368};
  assign T368 = T369;
  assign T369 = T370 != 2'h0;
  assign T370 = T354[9:8];
  assign T371 = T372;
  assign T372 = T373 != 2'h0;
  assign T373 = T354[11:10];
  assign T374 = T375;
  assign T375 = T376 != 2'h0;
  assign T376 = T354[13:12];
  assign T377 = {T393, T378};
  assign T378 = {T386, T379};
  assign T379 = {T383, T380};
  assign T380 = T381;
  assign T381 = T382 != 2'h0;
  assign T382 = T354[15:14];
  assign T383 = T384;
  assign T384 = T385 != 2'h0;
  assign T385 = T354[17:16];
  assign T386 = {T390, T387};
  assign T387 = T388;
  assign T388 = T389 != 2'h0;
  assign T389 = T354[19:18];
  assign T390 = T391;
  assign T391 = T392 != 2'h0;
  assign T392 = T354[21:20];
  assign T393 = {T401, T394};
  assign T394 = {T398, T395};
  assign T395 = T396;
  assign T396 = T397 != 2'h0;
  assign T397 = T354[23:22];
  assign T398 = T399;
  assign T399 = T400 != 2'h0;
  assign T400 = T354[25:24];
  assign T401 = T402;
  assign T402 = T403 != 1'h0;
  assign T403 = T354[26];
  assign T404 = T405 != 3'h0;
  assign T405 = notCDom_mainSig[2:0];
  assign notCDom_mainSig = T406[109:52];
  assign T406 = notCDom_absSigSum << notCDom_nearNormDist;
  assign notCDom_nearNormDist = T562 << 1'h1;
  assign T407 = notCDom_mainSig >> 2'h3;
  assign CDom_sig = {T520, T408};
  assign T408 = T414 | CDom_absSigSumExtra;
  assign CDom_absSigSumExtra = io_fromPreMul_doSubMags ? T411 : T409;
  assign T409 = T410 != 54'h0;
  assign T410 = sigSum[54:1];
  assign T411 = T412 != 53'h0;
  assign T412 = ~ T413;
  assign T413 = sigSum[53:1];
  assign T414 = T517 | CDom_reduced4SigExtra;
  assign CDom_reduced4SigExtra = T415 != 14'h0;
  assign T415 = T453 & T683;
  assign T683 = {1'h0, T416};
  assign T416 = {T434, T417};
  assign T417 = {T424, T418};
  assign T418 = T419[4];
  assign T419 = T420[12:8];
  assign T420 = T421[13:1];
  assign T421 = $signed(17'h10000) >>> T422;
  assign T422 = ~ T423;
  assign T423 = io_fromPreMul_CDom_CAlignDist >> 2'h2;
  assign T424 = {T430, T425};
  assign T425 = {T429, T426};
  assign T426 = T427[1];
  assign T427 = T428[3:2];
  assign T428 = T419[3:0];
  assign T429 = T427[0];
  assign T430 = {T433, T431};
  assign T431 = T432[1];
  assign T432 = T428[1:0];
  assign T433 = T432[0];
  assign T434 = T451 | T435;
  assign T435 = T436 & 8'haa;
  assign T436 = T437 << 1'h1;
  assign T437 = T438[6:0];
  assign T438 = T449 | T439;
  assign T439 = T440 & 8'hcc;
  assign T440 = T441 << 2'h2;
  assign T441 = T442[5:0];
  assign T442 = T447 | T443;
  assign T443 = T444 & 8'hf0;
  assign T444 = T445 << 3'h4;
  assign T445 = T446[3:0];
  assign T446 = T420[7:0];
  assign T447 = T684 & 8'hf;
  assign T684 = {4'h0, T448};
  assign T448 = T446 >> 3'h4;
  assign T449 = T685 & 8'h33;
  assign T685 = {2'h0, T450};
  assign T450 = T442 >> 2'h2;
  assign T451 = T686 & 8'h55;
  assign T686 = {1'h0, T452};
  assign T452 = T438 >> 1'h1;
  assign T453 = T454;
  assign T454 = {T490, T455};
  assign T455 = {T479, T456};
  assign T456 = {T472, T457};
  assign T457 = {T469, T458};
  assign T458 = T459;
  assign T459 = T460 != 4'h0;
  assign T460 = T461[3:0];
  assign T461 = T462 << 2'h2;
  assign T462 = CDom_absSigSum[52:0];
  assign CDom_absSigSum = io_fromPreMul_doSubMags ? T467 : T463;
  assign T463 = {1'h0, T464};
  assign T464 = {T466, T465};
  assign T465 = sigSum[159:55];
  assign T466 = io_fromPreMul_highAlignedSigC[54:53];
  assign T467 = ~ T468;
  assign T468 = sigSum[161:54];
  assign T469 = T470;
  assign T470 = T471 != 4'h0;
  assign T471 = T461[7:4];
  assign T472 = {T476, T473};
  assign T473 = T474;
  assign T474 = T475 != 4'h0;
  assign T475 = T461[11:8];
  assign T476 = T477;
  assign T477 = T478 != 4'h0;
  assign T478 = T461[15:12];
  assign T479 = {T487, T480};
  assign T480 = {T484, T481};
  assign T481 = T482;
  assign T482 = T483 != 4'h0;
  assign T483 = T461[19:16];
  assign T484 = T485;
  assign T485 = T486 != 4'h0;
  assign T486 = T461[23:20];
  assign T487 = T488;
  assign T488 = T489 != 4'h0;
  assign T489 = T461[27:24];
  assign T490 = {T506, T491};
  assign T491 = {T499, T492};
  assign T492 = {T496, T493};
  assign T493 = T494;
  assign T494 = T495 != 4'h0;
  assign T495 = T461[31:28];
  assign T496 = T497;
  assign T497 = T498 != 4'h0;
  assign T498 = T461[35:32];
  assign T499 = {T503, T500};
  assign T500 = T501;
  assign T501 = T502 != 4'h0;
  assign T502 = T461[39:36];
  assign T503 = T504;
  assign T504 = T505 != 4'h0;
  assign T505 = T461[43:40];
  assign T506 = {T514, T507};
  assign T507 = {T511, T508};
  assign T508 = T509;
  assign T509 = T510 != 4'h0;
  assign T510 = T461[47:44];
  assign T511 = T512;
  assign T512 = T513 != 4'h0;
  assign T513 = T461[51:48];
  assign T514 = T515;
  assign T515 = T516 != 3'h0;
  assign T516 = T461[54:52];
  assign T517 = T518 != 3'h0;
  assign T518 = CDom_mainSig[2:0];
  assign CDom_mainSig = T519[107:50];
  assign T519 = CDom_absSigSum << io_fromPreMul_CDom_CAlignDist;
  assign T520 = CDom_mainSig >> 2'h3;
  assign io_rawOut_sExp = T521;
  assign T521 = io_fromPreMul_CIsDominant ? CDom_sExp : notCDom_sExp;
  assign notCDom_sExp = io_fromPreMul_sExpSum - T687;
  assign T687 = {T688, T522};
  assign T522 = T523;
  assign T523 = {1'h0, notCDom_nearNormDist};
  assign T688 = T689 ? 5'h1f : 5'h0;
  assign T689 = T522[7];
  assign CDom_sExp = io_fromPreMul_sExpSum - T690;
  assign T690 = {T691, T524};
  assign T524 = T525;
  assign T525 = {1'h0, io_fromPreMul_doSubMags};
  assign T691 = T692 ? 11'h7ff : 11'h0;
  assign T692 = T524[1];
  assign io_rawOut_sign = T526;
  assign T526 = T535 | T527;
  assign T527 = T531 & T528;
  assign T528 = io_fromPreMul_CIsDominant ? CDom_sign : notCDom_sign;
  assign notCDom_sign = notCDom_completeCancellation ? roundingMode_min : T529;
  assign T529 = io_fromPreMul_signProd ^ notCDom_signSigSum;
  assign roundingMode_min = io_roundingMode == 3'h2;
  assign notCDom_completeCancellation = T530 == 2'h0;
  assign T530 = notCDom_sig[55:54];
  assign CDom_sign = io_fromPreMul_signProd ^ io_fromPreMul_doSubMags;
  assign T531 = T534 & T532;
  assign T532 = notNaN_addZeros ^ 1'h1;
  assign notNaN_addZeros = T533 & io_fromPreMul_isZeroC;
  assign T533 = io_fromPreMul_isZeroA | io_fromPreMul_isZeroB;
  assign T534 = notNaN_isInfOut ^ 1'h1;
  assign notNaN_isInfOut = notNaN_isInfProd | io_fromPreMul_isInfC;
  assign notNaN_isInfProd = io_fromPreMul_isInfA | io_fromPreMul_isInfB;
  assign T535 = T539 | T536;
  assign T536 = T538 & T537;
  assign T537 = io_fromPreMul_signProd | CDom_sign;
  assign T538 = notNaN_addZeros & roundingMode_min;
  assign T539 = T544 | T540;
  assign T540 = T541 & CDom_sign;
  assign T541 = T542 & io_fromPreMul_signProd;
  assign T542 = notNaN_addZeros & T543;
  assign T543 = roundingMode_min ^ 1'h1;
  assign T544 = T546 | T545;
  assign T545 = io_fromPreMul_isInfC & CDom_sign;
  assign T546 = notNaN_isInfProd & io_fromPreMul_signProd;
  assign io_rawOut_isZero = T547;
  assign T547 = notNaN_addZeros | T548;
  assign T548 = T549 & notCDom_completeCancellation;
  assign T549 = io_fromPreMul_CIsDominant ^ 1'h1;
  assign io_rawOut_isInf = notNaN_isInfOut;
  assign io_rawOut_isNaN = T550;
  assign T550 = io_fromPreMul_isNaNAOrB | io_fromPreMul_isNaNC;
  assign io_invalidExc = T551;
  assign T551 = T557 | T552;
  assign T552 = T553 & io_fromPreMul_doSubMags;
  assign T553 = T554 & io_fromPreMul_isInfC;
  assign T554 = T556 & T555;
  assign T555 = io_fromPreMul_isInfA | io_fromPreMul_isInfB;
  assign T556 = io_fromPreMul_isNaNAOrB ^ 1'h1;
  assign T557 = T559 | T558;
  assign T558 = io_fromPreMul_isZeroA & io_fromPreMul_isInfB;
  assign T559 = io_fromPreMul_isSigNaNAny | T560;
  assign T560 = io_fromPreMul_isInfA & io_fromPreMul_isZeroB;
endmodule

module RoundAnyRawFNToRecFN(
    input  io_invalidExc,
    input  io_infiniteExc,
    input  io_in_isNaN,
    input  io_in_isInf,
    input  io_in_isZero,
    input  io_in_sign,
    input [12:0] io_in_sExp,
    input [55:0] io_in_sig,
    input [2:0] io_roundingMode,
    input  io_detectTininess,
    output[64:0] io_out,
    output[4:0] io_exceptionFlags
);

  wire[4:0] T0;
  wire[2:0] T1;
  wire[1:0] T2;
  wire inexact;
  wire T3;
  wire common_inexact;
  wire T4;
  wire T5;
  wire T6;
  wire[55:0] T7;
  wire[55:0] T8;
  wire[54:0] T9;
  wire[55:0] T10;
  wire[53:0] T11;
  wire[53:0] T240;
  wire doShiftSigDown1;
  wire[53:0] T12;
  wire[53:0] T13;
  wire[53:0] T241;
  wire[2:0] T14;
  wire[2:0] T15;
  wire[2:0] T16;
  wire[2:0] T17;
  wire[2:0] T18;
  wire T19;
  wire[2:0] T20;
  wire[64:0] T21;
  wire[5:0] T22;
  wire[6:0] T23;
  wire[7:0] T24;
  wire[8:0] T25;
  wire[9:0] T26;
  wire[10:0] T27;
  wire[11:0] T28;
  wire[11:0] T29;
  wire[1:0] T30;
  wire T31;
  wire[1:0] T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire[53:0] T38;
  wire[50:0] T39;
  wire[50:0] T40;
  wire[50:0] T41;
  wire[50:0] T42;
  wire[50:0] T43;
  wire[50:0] T44;
  wire[50:0] T45;
  wire[50:0] T46;
  wire[50:0] T47;
  wire[50:0] T48;
  wire[50:0] T49;
  wire[50:0] T50;
  wire[50:0] T51;
  wire[18:0] T52;
  wire[2:0] T53;
  wire T54;
  wire[2:0] T55;
  wire[18:0] T56;
  wire[50:0] T57;
  wire[64:0] T58;
  wire[5:0] T59;
  wire[6:0] T60;
  wire[7:0] T61;
  wire[8:0] T62;
  wire[1:0] T63;
  wire T64;
  wire[1:0] T65;
  wire T66;
  wire[15:0] T67;
  wire[15:0] T68;
  wire[15:0] T69;
  wire[14:0] T70;
  wire[15:0] T71;
  wire[15:0] T72;
  wire[15:0] T73;
  wire[13:0] T74;
  wire[15:0] T75;
  wire[15:0] T76;
  wire[15:0] T77;
  wire[11:0] T78;
  wire[15:0] T79;
  wire[15:0] T80;
  wire[15:0] T81;
  wire[7:0] T82;
  wire[15:0] T83;
  wire[15:0] T84;
  wire[15:0] T242;
  wire[7:0] T85;
  wire[15:0] T86;
  wire[15:0] T243;
  wire[11:0] T87;
  wire[15:0] T88;
  wire[15:0] T244;
  wire[13:0] T89;
  wire[15:0] T90;
  wire[15:0] T245;
  wire[14:0] T91;
  wire[31:0] T92;
  wire[31:0] T93;
  wire[31:0] T94;
  wire[30:0] T95;
  wire[31:0] T96;
  wire[31:0] T97;
  wire[31:0] T98;
  wire[29:0] T99;
  wire[31:0] T100;
  wire[31:0] T101;
  wire[31:0] T102;
  wire[27:0] T103;
  wire[31:0] T104;
  wire[31:0] T105;
  wire[31:0] T106;
  wire[23:0] T107;
  wire[31:0] T108;
  wire[31:0] T109;
  wire[31:0] T110;
  wire[15:0] T111;
  wire[31:0] T112;
  wire[31:0] T113;
  wire[31:0] T246;
  wire[15:0] T114;
  wire[31:0] T115;
  wire[31:0] T247;
  wire[23:0] T116;
  wire[31:0] T117;
  wire[31:0] T248;
  wire[27:0] T118;
  wire[31:0] T119;
  wire[31:0] T249;
  wire[29:0] T120;
  wire[31:0] T121;
  wire[31:0] T250;
  wire[30:0] T122;
  wire T123;
  wire T124;
  wire T125;
  wire T126;
  wire T127;
  wire T128;
  wire[55:0] adjustedSig;
  wire T129;
  wire[55:0] T130;
  wire[55:0] T131;
  wire[55:0] T132;
  wire common_totalUnderflow;
  wire T133;
  wire[15:0] T134;
  wire[14:0] T251;
  wire[3:0] T135;
  wire[3:0] T136;
  wire[2:0] T137;
  wire[55:0] T138;
  wire[54:0] T139;
  wire[54:0] T140;
  wire[54:0] T141;
  wire T142;
  wire roundingMode_odd;
  wire[54:0] T252;
  wire[53:0] T143;
  wire[55:0] T144;
  wire[55:0] T145;
  wire[55:0] T146;
  wire[54:0] T147;
  wire[54:0] T148;
  wire[54:0] T149;
  wire T150;
  wire T151;
  wire T152;
  wire roundingMode_near_even;
  wire[55:0] T153;
  wire[54:0] T253;
  wire[53:0] T154;
  wire[55:0] T155;
  wire T156;
  wire T157;
  wire roundMagUp;
  wire T158;
  wire T159;
  wire roundingMode_max;
  wire T160;
  wire roundingMode_min;
  wire T161;
  wire T162;
  wire roundingMode_near_maxMag;
  wire[10:0] T254;
  wire T255;
  wire[13:0] T256;
  wire T257;
  wire commonCase;
  wire T163;
  wire T164;
  wire T165;
  wire notNaN_isSpecialInfOut;
  wire T166;
  wire isNaNOut;
  wire underflow;
  wire common_underflow;
  wire T167;
  wire T168;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire T173;
  wire T174;
  wire[1:0] T175;
  wire T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  wire T182;
  wire T183;
  wire T184;
  wire T185;
  wire T186;
  wire T187;
  wire T188;
  wire T189;
  wire T190;
  wire T191;
  wire T192;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  wire T198;
  wire T199;
  wire[1:0] T200;
  wire overflow;
  wire common_overflow;
  wire T201;
  wire[5:0] T202;
  wire[1:0] T203;
  wire[64:0] T204;
  wire[63:0] T205;
  wire[51:0] fractOut;
  wire[51:0] T206;
  wire[51:0] T258;
  wire pegMaxFiniteMagOut;
  wire T207;
  wire overflow_roundMagUp;
  wire T208;
  wire[51:0] T209;
  wire[51:0] common_fractOut;
  wire[51:0] T210;
  wire[51:0] T211;
  wire[51:0] T212;
  wire[51:0] T213;
  wire T214;
  wire T215;
  wire[11:0] expOut;
  wire[11:0] T216;
  wire[11:0] T217;
  wire[11:0] T218;
  wire notNaN_isInfOut;
  wire T219;
  wire[11:0] T220;
  wire[11:0] T221;
  wire[11:0] T222;
  wire[11:0] T223;
  wire pegMinNonzeroMagOut;
  wire T224;
  wire T225;
  wire[11:0] T226;
  wire[11:0] T227;
  wire[11:0] T228;
  wire[11:0] T229;
  wire[11:0] T230;
  wire[11:0] T231;
  wire[11:0] T232;
  wire[11:0] T233;
  wire[11:0] T234;
  wire[11:0] T235;
  wire[11:0] T236;
  wire[11:0] T237;
  wire T238;
  wire[11:0] common_expOut;
  wire[11:0] T239;
  wire signOut;


  assign io_exceptionFlags = T0;
  assign T0 = {T203, T1};
  assign T1 = {overflow, T2};
  assign T2 = {underflow, inexact};
  assign inexact = overflow | T3;
  assign T3 = commonCase & common_inexact;
  assign common_inexact = T4;
  assign T4 = common_totalUnderflow | T5;
  assign T5 = T129 | T6;
  assign T6 = T7 != 56'h0;
  assign T7 = adjustedSig & T8;
  assign T8 = {1'h0, T9};
  assign T9 = T10 >> 1'h1;
  assign T10 = {T11, 2'h3};
  assign T11 = T12 | T240;
  assign T240 = {53'h0, doShiftSigDown1};
  assign doShiftSigDown1 = adjustedSig[55];
  assign T12 = T128 ? T13 : 54'h0;
  assign T13 = T127 ? T38 : T241;
  assign T241 = {51'h0, T14};
  assign T14 = T37 ? T15 : 3'h0;
  assign T15 = T36 ? T16 : 3'h0;
  assign T16 = T35 ? T17 : 3'h0;
  assign T17 = T34 ? T18 : 3'h0;
  assign T18 = {T30, T19};
  assign T19 = T20[2];
  assign T20 = T21[2:0];
  assign T21 = $signed(65'h10000000000000000) >>> T22;
  assign T22 = T23[5:0];
  assign T23 = T24[6:0];
  assign T24 = T25[7:0];
  assign T25 = T26[8:0];
  assign T26 = T27[9:0];
  assign T27 = T28[10:0];
  assign T28 = ~ T29;
  assign T29 = io_in_sExp[11:0];
  assign T30 = {T33, T31};
  assign T31 = T32[1];
  assign T32 = T20[1:0];
  assign T33 = T32[0];
  assign T34 = T23[6];
  assign T35 = T24[7];
  assign T36 = T25[8];
  assign T37 = T26[9];
  assign T38 = {T39, 3'h7};
  assign T39 = ~ T40;
  assign T40 = T126 ? 51'h0 : T41;
  assign T41 = ~ T42;
  assign T42 = ~ T43;
  assign T43 = T125 ? 51'h0 : T44;
  assign T44 = ~ T45;
  assign T45 = ~ T46;
  assign T46 = T124 ? 51'h0 : T47;
  assign T47 = ~ T48;
  assign T48 = ~ T49;
  assign T49 = T123 ? 51'h0 : T50;
  assign T50 = ~ T51;
  assign T51 = {T92, T52};
  assign T52 = {T67, T53};
  assign T53 = {T63, T54};
  assign T54 = T55[2];
  assign T55 = T56[18:16];
  assign T56 = T57[50:32];
  assign T57 = T58[63:13];
  assign T58 = $signed(65'h10000000000000000) >>> T59;
  assign T59 = T60[5:0];
  assign T60 = T61[6:0];
  assign T61 = T62[7:0];
  assign T62 = T26[8:0];
  assign T63 = {T66, T64};
  assign T64 = T65[1];
  assign T65 = T55[1:0];
  assign T66 = T65[0];
  assign T67 = T90 | T68;
  assign T68 = T69 & 16'haaaa;
  assign T69 = T70 << 1'h1;
  assign T70 = T71[14:0];
  assign T71 = T88 | T72;
  assign T72 = T73 & 16'hcccc;
  assign T73 = T74 << 2'h2;
  assign T74 = T75[13:0];
  assign T75 = T86 | T76;
  assign T76 = T77 & 16'hf0f0;
  assign T77 = T78 << 3'h4;
  assign T78 = T79[11:0];
  assign T79 = T84 | T80;
  assign T80 = T81 & 16'hff00;
  assign T81 = T82 << 4'h8;
  assign T82 = T83[7:0];
  assign T83 = T56[15:0];
  assign T84 = T242 & 16'hff;
  assign T242 = {8'h0, T85};
  assign T85 = T83 >> 4'h8;
  assign T86 = T243 & 16'hf0f;
  assign T243 = {4'h0, T87};
  assign T87 = T79 >> 3'h4;
  assign T88 = T244 & 16'h3333;
  assign T244 = {2'h0, T89};
  assign T89 = T75 >> 2'h2;
  assign T90 = T245 & 16'h5555;
  assign T245 = {1'h0, T91};
  assign T91 = T71 >> 1'h1;
  assign T92 = T121 | T93;
  assign T93 = T94 & 32'haaaaaaaa;
  assign T94 = T95 << 1'h1;
  assign T95 = T96[30:0];
  assign T96 = T119 | T97;
  assign T97 = T98 & 32'hcccccccc;
  assign T98 = T99 << 2'h2;
  assign T99 = T100[29:0];
  assign T100 = T117 | T101;
  assign T101 = T102 & 32'hf0f0f0f0;
  assign T102 = T103 << 3'h4;
  assign T103 = T104[27:0];
  assign T104 = T115 | T105;
  assign T105 = T106 & 32'hff00ff00;
  assign T106 = T107 << 4'h8;
  assign T107 = T108[23:0];
  assign T108 = T113 | T109;
  assign T109 = T110 & 32'hffff0000;
  assign T110 = T111 << 5'h10;
  assign T111 = T112[15:0];
  assign T112 = T57[31:0];
  assign T113 = T246 & 32'hffff;
  assign T246 = {16'h0, T114};
  assign T114 = T112 >> 5'h10;
  assign T115 = T247 & 32'hff00ff;
  assign T247 = {8'h0, T116};
  assign T116 = T108 >> 4'h8;
  assign T117 = T248 & 32'hf0f0f0f;
  assign T248 = {4'h0, T118};
  assign T118 = T104 >> 3'h4;
  assign T119 = T249 & 32'h33333333;
  assign T249 = {2'h0, T120};
  assign T120 = T100 >> 2'h2;
  assign T121 = T250 & 32'h55555555;
  assign T250 = {1'h0, T122};
  assign T122 = T96 >> 1'h1;
  assign T123 = T60[6];
  assign T124 = T61[7];
  assign T125 = T62[8];
  assign T126 = T26[9];
  assign T127 = T27[10];
  assign T128 = T28[11];
  assign adjustedSig = io_in_sig << 1'h0;
  assign T129 = T130 != 56'h0;
  assign T130 = adjustedSig & T131;
  assign T131 = T132 & T10;
  assign T132 = ~ T8;
  assign common_totalUnderflow = T133;
  assign T133 = $signed(T134) < $signed(11'h3ce);
  assign T134 = T256 + T251;
  assign T251 = {T254, T135};
  assign T135 = T136;
  assign T136 = {1'h0, T137};
  assign T137 = T138 >> 6'h35;
  assign T138 = T156 ? T146 : T139;
  assign T139 = T252 | T140;
  assign T140 = T142 ? T141 : 55'h0;
  assign T141 = T131 >> 1'h1;
  assign T142 = roundingMode_odd & T5;
  assign roundingMode_odd = io_roundingMode == 3'h6;
  assign T252 = {1'h0, T143};
  assign T143 = T144 >> 2'h2;
  assign T144 = adjustedSig & T145;
  assign T145 = ~ T10;
  assign T146 = T153 & T147;
  assign T147 = ~ T148;
  assign T148 = T150 ? T149 : 55'h0;
  assign T149 = T10 >> 1'h1;
  assign T150 = T152 & T151;
  assign T151 = T6 ^ 1'h1;
  assign T152 = roundingMode_near_even & T129;
  assign roundingMode_near_even = io_roundingMode == 3'h0;
  assign T153 = T253 + 55'h1;
  assign T253 = {1'h0, T154};
  assign T154 = T155 >> 2'h2;
  assign T155 = adjustedSig | T10;
  assign T156 = T161 | T157;
  assign T157 = roundMagUp & T5;
  assign roundMagUp = T160 | T158;
  assign T158 = roundingMode_max & T159;
  assign T159 = io_in_sign ^ 1'h1;
  assign roundingMode_max = io_roundingMode == 3'h3;
  assign T160 = roundingMode_min & io_in_sign;
  assign roundingMode_min = io_roundingMode == 3'h2;
  assign T161 = T162 & T129;
  assign T162 = roundingMode_near_even | roundingMode_near_maxMag;
  assign roundingMode_near_maxMag = io_roundingMode == 3'h4;
  assign T254 = T255 ? 11'h7ff : 11'h0;
  assign T255 = T135[2];
  assign T256 = {T257, io_in_sExp};
  assign T257 = io_in_sExp[12];
  assign commonCase = T164 & T163;
  assign T163 = io_in_isZero ^ 1'h1;
  assign T164 = T166 & T165;
  assign T165 = notNaN_isSpecialInfOut ^ 1'h1;
  assign notNaN_isSpecialInfOut = io_infiniteExc | io_in_isInf;
  assign T166 = isNaNOut ^ 1'h1;
  assign isNaNOut = io_invalidExc | io_in_isNaN;
  assign underflow = commonCase & common_underflow;
  assign common_underflow = T167;
  assign T167 = common_totalUnderflow | T168;
  assign T168 = T194 & T169;
  assign T169 = T170 ^ 1'h1;
  assign T170 = T183 & T171;
  assign T171 = T178 | T172;
  assign T172 = roundMagUp & T173;
  assign T173 = T176 | T174;
  assign T174 = T175 != 2'h0;
  assign T175 = adjustedSig[1:0];
  assign T176 = doShiftSigDown1 & T177;
  assign T177 = adjustedSig[2];
  assign T178 = T182 & T179;
  assign T179 = doShiftSigDown1 ? T181 : T180;
  assign T180 = adjustedSig[1];
  assign T181 = adjustedSig[2];
  assign T182 = roundingMode_near_even | roundingMode_near_maxMag;
  assign T183 = T184 & T129;
  assign T184 = T188 & T185;
  assign T185 = doShiftSigDown1 ? T187 : T186;
  assign T186 = T138[53];
  assign T187 = T138[54];
  assign T188 = T193 & T189;
  assign T189 = T190 ^ 1'h1;
  assign T190 = doShiftSigDown1 ? T192 : T191;
  assign T191 = T10[3];
  assign T192 = T10[4];
  assign T193 = io_detectTininess == 1'h1;
  assign T194 = T198 & T195;
  assign T195 = doShiftSigDown1 ? T197 : T196;
  assign T196 = T10[2];
  assign T197 = T10[3];
  assign T198 = T5 & T199;
  assign T199 = $signed(T200) <= $signed(1'h0);
  assign T200 = $signed(io_in_sExp) >>> 4'hb;
  assign overflow = commonCase & common_overflow;
  assign common_overflow = T201;
  assign T201 = $signed(3'h3) <= $signed(T202);
  assign T202 = $signed(T134) >>> 4'ha;
  assign T203 = {io_invalidExc, io_infiniteExc};
  assign io_out = T204;
  assign T204 = {signOut, T205};
  assign T205 = {expOut, fractOut};
  assign fractOut = T209 | T206;
  assign T206 = 52'h0 - T258;
  assign T258 = {51'h0, pegMaxFiniteMagOut};
  assign pegMaxFiniteMagOut = overflow & T207;
  assign T207 = overflow_roundMagUp ^ 1'h1;
  assign overflow_roundMagUp = T208 | roundMagUp;
  assign T208 = roundingMode_near_even | roundingMode_near_maxMag;
  assign T209 = T214 ? T213 : common_fractOut;
  assign common_fractOut = T210;
  assign T210 = doShiftSigDown1 ? T212 : T211;
  assign T211 = T138[51:0];
  assign T212 = T138[52:1];
  assign T213 = isNaNOut ? 52'h8000000000000 : 52'h0;
  assign T214 = T215 | common_totalUnderflow;
  assign T215 = isNaNOut | io_in_isZero;
  assign expOut = T217 | T216;
  assign T216 = isNaNOut ? 12'he00 : 12'h0;
  assign T217 = T220 | T218;
  assign T218 = notNaN_isInfOut ? 12'hc00 : 12'h0;
  assign notNaN_isInfOut = notNaN_isSpecialInfOut | T219;
  assign T219 = overflow & overflow_roundMagUp;
  assign T220 = T222 | T221;
  assign T221 = pegMaxFiniteMagOut ? 12'hbff : 12'h0;
  assign T222 = T226 | T223;
  assign T223 = pegMinNonzeroMagOut ? 12'h3ce : 12'h0;
  assign pegMinNonzeroMagOut = T225 & T224;
  assign T224 = roundMagUp | roundingMode_odd;
  assign T225 = commonCase & common_totalUnderflow;
  assign T226 = T229 & T227;
  assign T227 = ~ T228;
  assign T228 = notNaN_isInfOut ? 12'h200 : 12'h0;
  assign T229 = T232 & T230;
  assign T230 = ~ T231;
  assign T231 = pegMaxFiniteMagOut ? 12'h400 : 12'h0;
  assign T232 = T235 & T233;
  assign T233 = ~ T234;
  assign T234 = pegMinNonzeroMagOut ? 12'hc31 : 12'h0;
  assign T235 = common_expOut & T236;
  assign T236 = ~ T237;
  assign T237 = T238 ? 12'he00 : 12'h0;
  assign T238 = io_in_isZero | common_totalUnderflow;
  assign common_expOut = T239;
  assign T239 = T134[11:0];
  assign signOut = isNaNOut ? 1'h0 : io_in_sign;
endmodule

module RoundRawFNToRecFN(
    input  io_invalidExc,
    input  io_infiniteExc,
    input  io_in_isNaN,
    input  io_in_isInf,
    input  io_in_isZero,
    input  io_in_sign,
    input [12:0] io_in_sExp,
    input [55:0] io_in_sig,
    input [2:0] io_roundingMode,
    input  io_detectTininess,
    output[64:0] io_out,
    output[4:0] io_exceptionFlags
);

  wire[64:0] roundAnyRawFNToRecFN_io_out;
  wire[4:0] roundAnyRawFNToRecFN_io_exceptionFlags;


  assign io_exceptionFlags = roundAnyRawFNToRecFN_io_exceptionFlags;
  assign io_out = roundAnyRawFNToRecFN_io_out;
  RoundAnyRawFNToRecFN roundAnyRawFNToRecFN(
       .io_invalidExc( io_invalidExc ),
       .io_infiniteExc( io_infiniteExc ),
       .io_in_isNaN( io_in_isNaN ),
       .io_in_isInf( io_in_isInf ),
       .io_in_isZero( io_in_isZero ),
       .io_in_sign( io_in_sign ),
       .io_in_sExp( io_in_sExp ),
       .io_in_sig( io_in_sig ),
       .io_roundingMode( io_roundingMode ),
       .io_detectTininess( io_detectTininess ),
       .io_out( roundAnyRawFNToRecFN_io_out ),
       .io_exceptionFlags( roundAnyRawFNToRecFN_io_exceptionFlags )
  );
endmodule

module MulAddRecFN(
    input [1:0] io_op,
    input [64:0] io_a,
    input [64:0] io_b,
    input [64:0] io_c,
    input [2:0] io_roundingMode,
    input  io_detectTininess,
    output[64:0] io_out,
    output[4:0] io_exceptionFlags
);

  wire[106:0] mulAddResult;
  wire[106:0] T1;
  wire[106:0] T2;
  wire[105:0] T0;
  wire[52:0] mulAddRecFNToRaw_preMul_io_mulAddA;
  wire[52:0] mulAddRecFNToRaw_preMul_io_mulAddB;
  wire[105:0] mulAddRecFNToRaw_preMul_io_mulAddC;
  wire mulAddRecFNToRaw_preMul_io_toPostMul_isSigNaNAny;
  wire mulAddRecFNToRaw_preMul_io_toPostMul_isNaNAOrB;
  wire mulAddRecFNToRaw_preMul_io_toPostMul_isInfA;
  wire mulAddRecFNToRaw_preMul_io_toPostMul_isZeroA;
  wire mulAddRecFNToRaw_preMul_io_toPostMul_isInfB;
  wire mulAddRecFNToRaw_preMul_io_toPostMul_isZeroB;
  wire mulAddRecFNToRaw_preMul_io_toPostMul_signProd;
  wire mulAddRecFNToRaw_preMul_io_toPostMul_isNaNC;
  wire mulAddRecFNToRaw_preMul_io_toPostMul_isInfC;
  wire mulAddRecFNToRaw_preMul_io_toPostMul_isZeroC;
  wire[12:0] mulAddRecFNToRaw_preMul_io_toPostMul_sExpSum;
  wire mulAddRecFNToRaw_preMul_io_toPostMul_doSubMags;
  wire mulAddRecFNToRaw_preMul_io_toPostMul_CIsDominant;
  wire[5:0] mulAddRecFNToRaw_preMul_io_toPostMul_CDom_CAlignDist;
  wire[54:0] mulAddRecFNToRaw_preMul_io_toPostMul_highAlignedSigC;
  wire mulAddRecFNToRaw_preMul_io_toPostMul_bit0AlignedSigC;
  wire mulAddRecFNToRaw_postMul_io_invalidExc;
  wire mulAddRecFNToRaw_postMul_io_rawOut_isNaN;
  wire mulAddRecFNToRaw_postMul_io_rawOut_isInf;
  wire mulAddRecFNToRaw_postMul_io_rawOut_isZero;
  wire mulAddRecFNToRaw_postMul_io_rawOut_sign;
  wire[12:0] mulAddRecFNToRaw_postMul_io_rawOut_sExp;
  wire[55:0] mulAddRecFNToRaw_postMul_io_rawOut_sig;
  wire[64:0] roundRawFNToRecFN_io_out;
  wire[4:0] roundRawFNToRecFN_io_exceptionFlags;


  assign mulAddResult = T2 + T1;
  assign T1 = {1'h0, mulAddRecFNToRaw_preMul_io_mulAddC};
  assign T2 = {1'h0, T0};
  assign T0 = mulAddRecFNToRaw_preMul_io_mulAddA * mulAddRecFNToRaw_preMul_io_mulAddB;
  assign io_exceptionFlags = roundRawFNToRecFN_io_exceptionFlags;
  assign io_out = roundRawFNToRecFN_io_out;
  MulAddRecFNToRaw_preMul mulAddRecFNToRaw_preMul(
       .io_op( io_op ),
       .io_a( io_a ),
       .io_b( io_b ),
       .io_c( io_c ),
       .io_mulAddA( mulAddRecFNToRaw_preMul_io_mulAddA ),
       .io_mulAddB( mulAddRecFNToRaw_preMul_io_mulAddB ),
       .io_mulAddC( mulAddRecFNToRaw_preMul_io_mulAddC ),
       .io_toPostMul_isSigNaNAny( mulAddRecFNToRaw_preMul_io_toPostMul_isSigNaNAny ),
       .io_toPostMul_isNaNAOrB( mulAddRecFNToRaw_preMul_io_toPostMul_isNaNAOrB ),
       .io_toPostMul_isInfA( mulAddRecFNToRaw_preMul_io_toPostMul_isInfA ),
       .io_toPostMul_isZeroA( mulAddRecFNToRaw_preMul_io_toPostMul_isZeroA ),
       .io_toPostMul_isInfB( mulAddRecFNToRaw_preMul_io_toPostMul_isInfB ),
       .io_toPostMul_isZeroB( mulAddRecFNToRaw_preMul_io_toPostMul_isZeroB ),
       .io_toPostMul_signProd( mulAddRecFNToRaw_preMul_io_toPostMul_signProd ),
       .io_toPostMul_isNaNC( mulAddRecFNToRaw_preMul_io_toPostMul_isNaNC ),
       .io_toPostMul_isInfC( mulAddRecFNToRaw_preMul_io_toPostMul_isInfC ),
       .io_toPostMul_isZeroC( mulAddRecFNToRaw_preMul_io_toPostMul_isZeroC ),
       .io_toPostMul_sExpSum( mulAddRecFNToRaw_preMul_io_toPostMul_sExpSum ),
       .io_toPostMul_doSubMags( mulAddRecFNToRaw_preMul_io_toPostMul_doSubMags ),
       .io_toPostMul_CIsDominant( mulAddRecFNToRaw_preMul_io_toPostMul_CIsDominant ),
       .io_toPostMul_CDom_CAlignDist( mulAddRecFNToRaw_preMul_io_toPostMul_CDom_CAlignDist ),
       .io_toPostMul_highAlignedSigC( mulAddRecFNToRaw_preMul_io_toPostMul_highAlignedSigC ),
       .io_toPostMul_bit0AlignedSigC( mulAddRecFNToRaw_preMul_io_toPostMul_bit0AlignedSigC )
  );
  MulAddRecFNToRaw_postMul mulAddRecFNToRaw_postMul(
       .io_fromPreMul_isSigNaNAny( mulAddRecFNToRaw_preMul_io_toPostMul_isSigNaNAny ),
       .io_fromPreMul_isNaNAOrB( mulAddRecFNToRaw_preMul_io_toPostMul_isNaNAOrB ),
       .io_fromPreMul_isInfA( mulAddRecFNToRaw_preMul_io_toPostMul_isInfA ),
       .io_fromPreMul_isZeroA( mulAddRecFNToRaw_preMul_io_toPostMul_isZeroA ),
       .io_fromPreMul_isInfB( mulAddRecFNToRaw_preMul_io_toPostMul_isInfB ),
       .io_fromPreMul_isZeroB( mulAddRecFNToRaw_preMul_io_toPostMul_isZeroB ),
       .io_fromPreMul_signProd( mulAddRecFNToRaw_preMul_io_toPostMul_signProd ),
       .io_fromPreMul_isNaNC( mulAddRecFNToRaw_preMul_io_toPostMul_isNaNC ),
       .io_fromPreMul_isInfC( mulAddRecFNToRaw_preMul_io_toPostMul_isInfC ),
       .io_fromPreMul_isZeroC( mulAddRecFNToRaw_preMul_io_toPostMul_isZeroC ),
       .io_fromPreMul_sExpSum( mulAddRecFNToRaw_preMul_io_toPostMul_sExpSum ),
       .io_fromPreMul_doSubMags( mulAddRecFNToRaw_preMul_io_toPostMul_doSubMags ),
       .io_fromPreMul_CIsDominant( mulAddRecFNToRaw_preMul_io_toPostMul_CIsDominant ),
       .io_fromPreMul_CDom_CAlignDist( mulAddRecFNToRaw_preMul_io_toPostMul_CDom_CAlignDist ),
       .io_fromPreMul_highAlignedSigC( mulAddRecFNToRaw_preMul_io_toPostMul_highAlignedSigC ),
       .io_fromPreMul_bit0AlignedSigC( mulAddRecFNToRaw_preMul_io_toPostMul_bit0AlignedSigC ),
       .io_mulAddResult( mulAddResult ),
       .io_roundingMode( io_roundingMode ),
       .io_invalidExc( mulAddRecFNToRaw_postMul_io_invalidExc ),
       .io_rawOut_isNaN( mulAddRecFNToRaw_postMul_io_rawOut_isNaN ),
       .io_rawOut_isInf( mulAddRecFNToRaw_postMul_io_rawOut_isInf ),
       .io_rawOut_isZero( mulAddRecFNToRaw_postMul_io_rawOut_isZero ),
       .io_rawOut_sign( mulAddRecFNToRaw_postMul_io_rawOut_sign ),
       .io_rawOut_sExp( mulAddRecFNToRaw_postMul_io_rawOut_sExp ),
       .io_rawOut_sig( mulAddRecFNToRaw_postMul_io_rawOut_sig )
  );
  RoundRawFNToRecFN roundRawFNToRecFN(
       .io_invalidExc( mulAddRecFNToRaw_postMul_io_invalidExc ),
       .io_infiniteExc( 1'h0 ),
       .io_in_isNaN( mulAddRecFNToRaw_postMul_io_rawOut_isNaN ),
       .io_in_isInf( mulAddRecFNToRaw_postMul_io_rawOut_isInf ),
       .io_in_isZero( mulAddRecFNToRaw_postMul_io_rawOut_isZero ),
       .io_in_sign( mulAddRecFNToRaw_postMul_io_rawOut_sign ),
       .io_in_sExp( mulAddRecFNToRaw_postMul_io_rawOut_sExp ),
       .io_in_sig( mulAddRecFNToRaw_postMul_io_rawOut_sig ),
       .io_roundingMode( io_roundingMode ),
       .io_detectTininess( io_detectTininess ),
       .io_out( roundRawFNToRecFN_io_out ),
       .io_exceptionFlags( roundRawFNToRecFN_io_exceptionFlags )
  );
endmodule

module ValExec_MulAddRecF64(
    input [63:0] io_a,
    input [63:0] io_b,
    input [63:0] io_c,
    input [2:0] io_roundingMode,
    input  io_detectTininess,
    input [63:0] io_expected_out,
    input [4:0] io_expected_exceptionFlags,
    output[64:0] io_expected_recOut,
    output[64:0] io_actual_out,
    output[4:0] io_actual_exceptionFlags,
    output io_check,
    output io_pass
);

  wire[64:0] T0;
  wire[60:0] T1;
  wire[51:0] T2;
  wire[53:0] T3;
  wire[53:0] T4;
  wire[52:0] T5;
  wire[51:0] T6;
  wire[51:0] T7;
  wire[51:0] T8;
  wire[50:0] T9;
  wire[114:0] T10;
  wire[5:0] T452;
  wire[5:0] T453;
  wire[5:0] T454;
  wire[5:0] T455;
  wire[5:0] T456;
  wire[5:0] T457;
  wire[5:0] T458;
  wire[5:0] T459;
  wire[5:0] T460;
  wire[5:0] T461;
  wire[5:0] T462;
  wire[5:0] T463;
  wire[5:0] T464;
  wire[5:0] T465;
  wire[5:0] T466;
  wire[5:0] T467;
  wire[5:0] T468;
  wire[5:0] T469;
  wire[5:0] T470;
  wire[5:0] T471;
  wire[5:0] T472;
  wire[5:0] T473;
  wire[5:0] T474;
  wire[5:0] T475;
  wire[5:0] T476;
  wire[5:0] T477;
  wire[5:0] T478;
  wire[5:0] T479;
  wire[5:0] T480;
  wire[5:0] T481;
  wire[5:0] T482;
  wire[5:0] T483;
  wire[5:0] T484;
  wire[5:0] T485;
  wire[5:0] T486;
  wire[5:0] T487;
  wire[5:0] T488;
  wire[5:0] T489;
  wire[5:0] T490;
  wire[5:0] T491;
  wire[5:0] T492;
  wire[5:0] T493;
  wire[5:0] T494;
  wire[5:0] T495;
  wire[5:0] T496;
  wire[5:0] T497;
  wire[5:0] T498;
  wire[5:0] T499;
  wire[5:0] T500;
  wire[5:0] T501;
  wire[5:0] T502;
  wire T503;
  wire[51:0] T12;
  wire[19:0] T13;
  wire[3:0] T14;
  wire[1:0] T15;
  wire T16;
  wire[1:0] T17;
  wire[3:0] T18;
  wire[19:0] T19;
  wire T20;
  wire[1:0] T21;
  wire T22;
  wire[1:0] T23;
  wire T24;
  wire[15:0] T25;
  wire[15:0] T26;
  wire[15:0] T27;
  wire[14:0] T28;
  wire[15:0] T29;
  wire[15:0] T30;
  wire[15:0] T31;
  wire[13:0] T32;
  wire[15:0] T33;
  wire[15:0] T34;
  wire[15:0] T35;
  wire[11:0] T36;
  wire[15:0] T37;
  wire[15:0] T38;
  wire[15:0] T39;
  wire[7:0] T40;
  wire[15:0] T41;
  wire[15:0] T42;
  wire[15:0] T504;
  wire[7:0] T43;
  wire[15:0] T44;
  wire[15:0] T505;
  wire[11:0] T45;
  wire[15:0] T46;
  wire[15:0] T506;
  wire[13:0] T47;
  wire[15:0] T48;
  wire[15:0] T507;
  wire[14:0] T49;
  wire[31:0] T50;
  wire[31:0] T51;
  wire[31:0] T52;
  wire[30:0] T53;
  wire[31:0] T54;
  wire[31:0] T55;
  wire[31:0] T56;
  wire[29:0] T57;
  wire[31:0] T58;
  wire[31:0] T59;
  wire[31:0] T60;
  wire[27:0] T61;
  wire[31:0] T62;
  wire[31:0] T63;
  wire[31:0] T64;
  wire[23:0] T65;
  wire[31:0] T66;
  wire[31:0] T67;
  wire[31:0] T68;
  wire[15:0] T69;
  wire[31:0] T70;
  wire[31:0] T71;
  wire[31:0] T508;
  wire[15:0] T72;
  wire[31:0] T73;
  wire[31:0] T509;
  wire[23:0] T74;
  wire[31:0] T75;
  wire[31:0] T510;
  wire[27:0] T76;
  wire[31:0] T77;
  wire[31:0] T511;
  wire[29:0] T78;
  wire[31:0] T79;
  wire[31:0] T512;
  wire[30:0] T80;
  wire T513;
  wire T514;
  wire T515;
  wire T516;
  wire T517;
  wire T518;
  wire T519;
  wire T520;
  wire T521;
  wire T522;
  wire T523;
  wire T524;
  wire T525;
  wire T526;
  wire T527;
  wire T528;
  wire T529;
  wire T530;
  wire T531;
  wire T532;
  wire T533;
  wire T534;
  wire T535;
  wire T536;
  wire T537;
  wire T538;
  wire T539;
  wire T540;
  wire T541;
  wire T542;
  wire T543;
  wire T544;
  wire T545;
  wire T546;
  wire T547;
  wire T548;
  wire T549;
  wire T550;
  wire T551;
  wire T552;
  wire T553;
  wire T554;
  wire T555;
  wire T556;
  wire T557;
  wire T558;
  wire T559;
  wire T560;
  wire T561;
  wire T562;
  wire T81;
  wire[10:0] T82;
  wire T83;
  wire T84;
  wire T85;
  wire[8:0] T86;
  wire[12:0] T87;
  wire[12:0] T88;
  wire[12:0] T89;
  wire[11:0] T90;
  wire[11:0] T91;
  wire[11:0] T563;
  wire[10:0] T92;
  wire[10:0] T564;
  wire[1:0] T93;
  wire[11:0] T94;
  wire[11:0] T565;
  wire[11:0] T95;
  wire[11:0] T566;
  wire[3:0] T96;
  wire[2:0] T97;
  wire[2:0] T567;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire[1:0] T102;
  wire[2:0] T103;
  wire[2:0] T104;
  wire T105;
  wire T106;
  wire T107;
  wire[64:0] T108;
  wire[60:0] T109;
  wire[51:0] T110;
  wire[53:0] T111;
  wire[53:0] T112;
  wire[52:0] T113;
  wire[51:0] T114;
  wire[51:0] T115;
  wire[51:0] T116;
  wire[50:0] T117;
  wire[114:0] T118;
  wire[5:0] T568;
  wire[5:0] T569;
  wire[5:0] T570;
  wire[5:0] T571;
  wire[5:0] T572;
  wire[5:0] T573;
  wire[5:0] T574;
  wire[5:0] T575;
  wire[5:0] T576;
  wire[5:0] T577;
  wire[5:0] T578;
  wire[5:0] T579;
  wire[5:0] T580;
  wire[5:0] T581;
  wire[5:0] T582;
  wire[5:0] T583;
  wire[5:0] T584;
  wire[5:0] T585;
  wire[5:0] T586;
  wire[5:0] T587;
  wire[5:0] T588;
  wire[5:0] T589;
  wire[5:0] T590;
  wire[5:0] T591;
  wire[5:0] T592;
  wire[5:0] T593;
  wire[5:0] T594;
  wire[5:0] T595;
  wire[5:0] T596;
  wire[5:0] T597;
  wire[5:0] T598;
  wire[5:0] T599;
  wire[5:0] T600;
  wire[5:0] T601;
  wire[5:0] T602;
  wire[5:0] T603;
  wire[5:0] T604;
  wire[5:0] T605;
  wire[5:0] T606;
  wire[5:0] T607;
  wire[5:0] T608;
  wire[5:0] T609;
  wire[5:0] T610;
  wire[5:0] T611;
  wire[5:0] T612;
  wire[5:0] T613;
  wire[5:0] T614;
  wire[5:0] T615;
  wire[5:0] T616;
  wire[5:0] T617;
  wire[5:0] T618;
  wire T619;
  wire[51:0] T120;
  wire[19:0] T121;
  wire[3:0] T122;
  wire[1:0] T123;
  wire T124;
  wire[1:0] T125;
  wire[3:0] T126;
  wire[19:0] T127;
  wire T128;
  wire[1:0] T129;
  wire T130;
  wire[1:0] T131;
  wire T132;
  wire[15:0] T133;
  wire[15:0] T134;
  wire[15:0] T135;
  wire[14:0] T136;
  wire[15:0] T137;
  wire[15:0] T138;
  wire[15:0] T139;
  wire[13:0] T140;
  wire[15:0] T141;
  wire[15:0] T142;
  wire[15:0] T143;
  wire[11:0] T144;
  wire[15:0] T145;
  wire[15:0] T146;
  wire[15:0] T147;
  wire[7:0] T148;
  wire[15:0] T149;
  wire[15:0] T150;
  wire[15:0] T620;
  wire[7:0] T151;
  wire[15:0] T152;
  wire[15:0] T621;
  wire[11:0] T153;
  wire[15:0] T154;
  wire[15:0] T622;
  wire[13:0] T155;
  wire[15:0] T156;
  wire[15:0] T623;
  wire[14:0] T157;
  wire[31:0] T158;
  wire[31:0] T159;
  wire[31:0] T160;
  wire[30:0] T161;
  wire[31:0] T162;
  wire[31:0] T163;
  wire[31:0] T164;
  wire[29:0] T165;
  wire[31:0] T166;
  wire[31:0] T167;
  wire[31:0] T168;
  wire[27:0] T169;
  wire[31:0] T170;
  wire[31:0] T171;
  wire[31:0] T172;
  wire[23:0] T173;
  wire[31:0] T174;
  wire[31:0] T175;
  wire[31:0] T176;
  wire[15:0] T177;
  wire[31:0] T178;
  wire[31:0] T179;
  wire[31:0] T624;
  wire[15:0] T180;
  wire[31:0] T181;
  wire[31:0] T625;
  wire[23:0] T182;
  wire[31:0] T183;
  wire[31:0] T626;
  wire[27:0] T184;
  wire[31:0] T185;
  wire[31:0] T627;
  wire[29:0] T186;
  wire[31:0] T187;
  wire[31:0] T628;
  wire[30:0] T188;
  wire T629;
  wire T630;
  wire T631;
  wire T632;
  wire T633;
  wire T634;
  wire T635;
  wire T636;
  wire T637;
  wire T638;
  wire T639;
  wire T640;
  wire T641;
  wire T642;
  wire T643;
  wire T644;
  wire T645;
  wire T646;
  wire T647;
  wire T648;
  wire T649;
  wire T650;
  wire T651;
  wire T652;
  wire T653;
  wire T654;
  wire T655;
  wire T656;
  wire T657;
  wire T658;
  wire T659;
  wire T660;
  wire T661;
  wire T662;
  wire T663;
  wire T664;
  wire T665;
  wire T666;
  wire T667;
  wire T668;
  wire T669;
  wire T670;
  wire T671;
  wire T672;
  wire T673;
  wire T674;
  wire T675;
  wire T676;
  wire T677;
  wire T678;
  wire T189;
  wire[10:0] T190;
  wire T191;
  wire T192;
  wire T193;
  wire[8:0] T194;
  wire[12:0] T195;
  wire[12:0] T196;
  wire[12:0] T197;
  wire[11:0] T198;
  wire[11:0] T199;
  wire[11:0] T679;
  wire[10:0] T200;
  wire[10:0] T680;
  wire[1:0] T201;
  wire[11:0] T202;
  wire[11:0] T681;
  wire[11:0] T203;
  wire[11:0] T682;
  wire[3:0] T204;
  wire[2:0] T205;
  wire[2:0] T683;
  wire T206;
  wire T207;
  wire T208;
  wire T209;
  wire[1:0] T210;
  wire[2:0] T211;
  wire[2:0] T212;
  wire T213;
  wire T214;
  wire T215;
  wire[64:0] T216;
  wire[60:0] T217;
  wire[51:0] T218;
  wire[53:0] T219;
  wire[53:0] T220;
  wire[52:0] T221;
  wire[51:0] T222;
  wire[51:0] T223;
  wire[51:0] T224;
  wire[50:0] T225;
  wire[114:0] T226;
  wire[5:0] T684;
  wire[5:0] T685;
  wire[5:0] T686;
  wire[5:0] T687;
  wire[5:0] T688;
  wire[5:0] T689;
  wire[5:0] T690;
  wire[5:0] T691;
  wire[5:0] T692;
  wire[5:0] T693;
  wire[5:0] T694;
  wire[5:0] T695;
  wire[5:0] T696;
  wire[5:0] T697;
  wire[5:0] T698;
  wire[5:0] T699;
  wire[5:0] T700;
  wire[5:0] T701;
  wire[5:0] T702;
  wire[5:0] T703;
  wire[5:0] T704;
  wire[5:0] T705;
  wire[5:0] T706;
  wire[5:0] T707;
  wire[5:0] T708;
  wire[5:0] T709;
  wire[5:0] T710;
  wire[5:0] T711;
  wire[5:0] T712;
  wire[5:0] T713;
  wire[5:0] T714;
  wire[5:0] T715;
  wire[5:0] T716;
  wire[5:0] T717;
  wire[5:0] T718;
  wire[5:0] T719;
  wire[5:0] T720;
  wire[5:0] T721;
  wire[5:0] T722;
  wire[5:0] T723;
  wire[5:0] T724;
  wire[5:0] T725;
  wire[5:0] T726;
  wire[5:0] T727;
  wire[5:0] T728;
  wire[5:0] T729;
  wire[5:0] T730;
  wire[5:0] T731;
  wire[5:0] T732;
  wire[5:0] T733;
  wire[5:0] T734;
  wire T735;
  wire[51:0] T228;
  wire[19:0] T229;
  wire[3:0] T230;
  wire[1:0] T231;
  wire T232;
  wire[1:0] T233;
  wire[3:0] T234;
  wire[19:0] T235;
  wire T236;
  wire[1:0] T237;
  wire T238;
  wire[1:0] T239;
  wire T240;
  wire[15:0] T241;
  wire[15:0] T242;
  wire[15:0] T243;
  wire[14:0] T244;
  wire[15:0] T245;
  wire[15:0] T246;
  wire[15:0] T247;
  wire[13:0] T248;
  wire[15:0] T249;
  wire[15:0] T250;
  wire[15:0] T251;
  wire[11:0] T252;
  wire[15:0] T253;
  wire[15:0] T254;
  wire[15:0] T255;
  wire[7:0] T256;
  wire[15:0] T257;
  wire[15:0] T258;
  wire[15:0] T736;
  wire[7:0] T259;
  wire[15:0] T260;
  wire[15:0] T737;
  wire[11:0] T261;
  wire[15:0] T262;
  wire[15:0] T738;
  wire[13:0] T263;
  wire[15:0] T264;
  wire[15:0] T739;
  wire[14:0] T265;
  wire[31:0] T266;
  wire[31:0] T267;
  wire[31:0] T268;
  wire[30:0] T269;
  wire[31:0] T270;
  wire[31:0] T271;
  wire[31:0] T272;
  wire[29:0] T273;
  wire[31:0] T274;
  wire[31:0] T275;
  wire[31:0] T276;
  wire[27:0] T277;
  wire[31:0] T278;
  wire[31:0] T279;
  wire[31:0] T280;
  wire[23:0] T281;
  wire[31:0] T282;
  wire[31:0] T283;
  wire[31:0] T284;
  wire[15:0] T285;
  wire[31:0] T286;
  wire[31:0] T287;
  wire[31:0] T740;
  wire[15:0] T288;
  wire[31:0] T289;
  wire[31:0] T741;
  wire[23:0] T290;
  wire[31:0] T291;
  wire[31:0] T742;
  wire[27:0] T292;
  wire[31:0] T293;
  wire[31:0] T743;
  wire[29:0] T294;
  wire[31:0] T295;
  wire[31:0] T744;
  wire[30:0] T296;
  wire T745;
  wire T746;
  wire T747;
  wire T748;
  wire T749;
  wire T750;
  wire T751;
  wire T752;
  wire T753;
  wire T754;
  wire T755;
  wire T756;
  wire T757;
  wire T758;
  wire T759;
  wire T760;
  wire T761;
  wire T762;
  wire T763;
  wire T764;
  wire T765;
  wire T766;
  wire T767;
  wire T768;
  wire T769;
  wire T770;
  wire T771;
  wire T772;
  wire T773;
  wire T774;
  wire T775;
  wire T776;
  wire T777;
  wire T778;
  wire T779;
  wire T780;
  wire T781;
  wire T782;
  wire T783;
  wire T784;
  wire T785;
  wire T786;
  wire T787;
  wire T788;
  wire T789;
  wire T790;
  wire T791;
  wire T792;
  wire T793;
  wire T794;
  wire T297;
  wire[10:0] T298;
  wire T299;
  wire T300;
  wire T301;
  wire[8:0] T302;
  wire[12:0] T303;
  wire[12:0] T304;
  wire[12:0] T305;
  wire[11:0] T306;
  wire[11:0] T307;
  wire[11:0] T795;
  wire[10:0] T308;
  wire[10:0] T796;
  wire[1:0] T309;
  wire[11:0] T310;
  wire[11:0] T797;
  wire[11:0] T311;
  wire[11:0] T798;
  wire[3:0] T312;
  wire[2:0] T313;
  wire[2:0] T799;
  wire T314;
  wire T315;
  wire T316;
  wire T317;
  wire[1:0] T318;
  wire[2:0] T319;
  wire[2:0] T320;
  wire T321;
  wire T322;
  wire T323;
  wire T324;
  wire T325;
  wire T326;
  wire T327;
  wire T328;
  wire T329;
  wire[3:0] T330;
  wire[3:0] T331;
  wire T332;
  wire[2:0] T333;
  wire T334;
  wire T335;
  wire[51:0] T336;
  wire[51:0] T337;
  wire T338;
  wire T339;
  wire T340;
  wire[2:0] T341;
  wire T342;
  wire[2:0] T343;
  wire[64:0] T344;
  wire[60:0] T345;
  wire[51:0] T346;
  wire[53:0] T347;
  wire[53:0] T348;
  wire[52:0] T349;
  wire[51:0] T350;
  wire[51:0] T351;
  wire[51:0] T352;
  wire[50:0] T353;
  wire[114:0] T354;
  wire[5:0] T800;
  wire[5:0] T801;
  wire[5:0] T802;
  wire[5:0] T803;
  wire[5:0] T804;
  wire[5:0] T805;
  wire[5:0] T806;
  wire[5:0] T807;
  wire[5:0] T808;
  wire[5:0] T809;
  wire[5:0] T810;
  wire[5:0] T811;
  wire[5:0] T812;
  wire[5:0] T813;
  wire[5:0] T814;
  wire[5:0] T815;
  wire[5:0] T816;
  wire[5:0] T817;
  wire[5:0] T818;
  wire[5:0] T819;
  wire[5:0] T820;
  wire[5:0] T821;
  wire[5:0] T822;
  wire[5:0] T823;
  wire[5:0] T824;
  wire[5:0] T825;
  wire[5:0] T826;
  wire[5:0] T827;
  wire[5:0] T828;
  wire[5:0] T829;
  wire[5:0] T830;
  wire[5:0] T831;
  wire[5:0] T832;
  wire[5:0] T833;
  wire[5:0] T834;
  wire[5:0] T835;
  wire[5:0] T836;
  wire[5:0] T837;
  wire[5:0] T838;
  wire[5:0] T839;
  wire[5:0] T840;
  wire[5:0] T841;
  wire[5:0] T842;
  wire[5:0] T843;
  wire[5:0] T844;
  wire[5:0] T845;
  wire[5:0] T846;
  wire[5:0] T847;
  wire[5:0] T848;
  wire[5:0] T849;
  wire[5:0] T850;
  wire T851;
  wire[51:0] T356;
  wire[19:0] T357;
  wire[3:0] T358;
  wire[1:0] T359;
  wire T360;
  wire[1:0] T361;
  wire[3:0] T362;
  wire[19:0] T363;
  wire T364;
  wire[1:0] T365;
  wire T366;
  wire[1:0] T367;
  wire T368;
  wire[15:0] T369;
  wire[15:0] T370;
  wire[15:0] T371;
  wire[14:0] T372;
  wire[15:0] T373;
  wire[15:0] T374;
  wire[15:0] T375;
  wire[13:0] T376;
  wire[15:0] T377;
  wire[15:0] T378;
  wire[15:0] T379;
  wire[11:0] T380;
  wire[15:0] T381;
  wire[15:0] T382;
  wire[15:0] T383;
  wire[7:0] T384;
  wire[15:0] T385;
  wire[15:0] T386;
  wire[15:0] T852;
  wire[7:0] T387;
  wire[15:0] T388;
  wire[15:0] T853;
  wire[11:0] T389;
  wire[15:0] T390;
  wire[15:0] T854;
  wire[13:0] T391;
  wire[15:0] T392;
  wire[15:0] T855;
  wire[14:0] T393;
  wire[31:0] T394;
  wire[31:0] T395;
  wire[31:0] T396;
  wire[30:0] T397;
  wire[31:0] T398;
  wire[31:0] T399;
  wire[31:0] T400;
  wire[29:0] T401;
  wire[31:0] T402;
  wire[31:0] T403;
  wire[31:0] T404;
  wire[27:0] T405;
  wire[31:0] T406;
  wire[31:0] T407;
  wire[31:0] T408;
  wire[23:0] T409;
  wire[31:0] T410;
  wire[31:0] T411;
  wire[31:0] T412;
  wire[15:0] T413;
  wire[31:0] T414;
  wire[31:0] T415;
  wire[31:0] T856;
  wire[15:0] T416;
  wire[31:0] T417;
  wire[31:0] T857;
  wire[23:0] T418;
  wire[31:0] T419;
  wire[31:0] T858;
  wire[27:0] T420;
  wire[31:0] T421;
  wire[31:0] T859;
  wire[29:0] T422;
  wire[31:0] T423;
  wire[31:0] T860;
  wire[30:0] T424;
  wire T861;
  wire T862;
  wire T863;
  wire T864;
  wire T865;
  wire T866;
  wire T867;
  wire T868;
  wire T869;
  wire T870;
  wire T871;
  wire T872;
  wire T873;
  wire T874;
  wire T875;
  wire T876;
  wire T877;
  wire T878;
  wire T879;
  wire T880;
  wire T881;
  wire T882;
  wire T883;
  wire T884;
  wire T885;
  wire T886;
  wire T887;
  wire T888;
  wire T889;
  wire T890;
  wire T891;
  wire T892;
  wire T893;
  wire T894;
  wire T895;
  wire T896;
  wire T897;
  wire T898;
  wire T899;
  wire T900;
  wire T901;
  wire T902;
  wire T903;
  wire T904;
  wire T905;
  wire T906;
  wire T907;
  wire T908;
  wire T909;
  wire T910;
  wire T425;
  wire[10:0] T426;
  wire T427;
  wire T428;
  wire T429;
  wire[8:0] T430;
  wire[12:0] T431;
  wire[12:0] T432;
  wire[12:0] T433;
  wire[11:0] T434;
  wire[11:0] T435;
  wire[11:0] T911;
  wire[10:0] T436;
  wire[10:0] T912;
  wire[1:0] T437;
  wire[11:0] T438;
  wire[11:0] T913;
  wire[11:0] T439;
  wire[11:0] T914;
  wire[3:0] T440;
  wire[2:0] T441;
  wire[2:0] T915;
  wire T442;
  wire T443;
  wire T444;
  wire T445;
  wire[1:0] T446;
  wire[2:0] T447;
  wire[2:0] T448;
  wire T449;
  wire T450;
  wire T451;
  wire[64:0] mulAddRecFN_io_out;
  wire[4:0] mulAddRecFN_io_exceptionFlags;


  assign T0 = {T96, T1};
  assign T1 = {T86, T2};
  assign T2 = T3[51:0];
  assign T3 = T4;
  assign T4 = {1'h0, T5};
  assign T5 = {T83, T6};
  assign T6 = T81 ? T8 : T7;
  assign T7 = io_c[51:0];
  assign T8 = T9 << 1'h1;
  assign T9 = T10[50:0];
  assign T10 = T7 << T452;
  assign T452 = T562 ? 1'h0 : T453;
  assign T453 = T561 ? 1'h1 : T454;
  assign T454 = T560 ? 2'h2 : T455;
  assign T455 = T559 ? 2'h3 : T456;
  assign T456 = T558 ? 3'h4 : T457;
  assign T457 = T557 ? 3'h5 : T458;
  assign T458 = T556 ? 3'h6 : T459;
  assign T459 = T555 ? 3'h7 : T460;
  assign T460 = T554 ? 4'h8 : T461;
  assign T461 = T553 ? 4'h9 : T462;
  assign T462 = T552 ? 4'ha : T463;
  assign T463 = T551 ? 4'hb : T464;
  assign T464 = T550 ? 4'hc : T465;
  assign T465 = T549 ? 4'hd : T466;
  assign T466 = T548 ? 4'he : T467;
  assign T467 = T547 ? 4'hf : T468;
  assign T468 = T546 ? 5'h10 : T469;
  assign T469 = T545 ? 5'h11 : T470;
  assign T470 = T544 ? 5'h12 : T471;
  assign T471 = T543 ? 5'h13 : T472;
  assign T472 = T542 ? 5'h14 : T473;
  assign T473 = T541 ? 5'h15 : T474;
  assign T474 = T540 ? 5'h16 : T475;
  assign T475 = T539 ? 5'h17 : T476;
  assign T476 = T538 ? 5'h18 : T477;
  assign T477 = T537 ? 5'h19 : T478;
  assign T478 = T536 ? 5'h1a : T479;
  assign T479 = T535 ? 5'h1b : T480;
  assign T480 = T534 ? 5'h1c : T481;
  assign T481 = T533 ? 5'h1d : T482;
  assign T482 = T532 ? 5'h1e : T483;
  assign T483 = T531 ? 5'h1f : T484;
  assign T484 = T530 ? 6'h20 : T485;
  assign T485 = T529 ? 6'h21 : T486;
  assign T486 = T528 ? 6'h22 : T487;
  assign T487 = T527 ? 6'h23 : T488;
  assign T488 = T526 ? 6'h24 : T489;
  assign T489 = T525 ? 6'h25 : T490;
  assign T490 = T524 ? 6'h26 : T491;
  assign T491 = T523 ? 6'h27 : T492;
  assign T492 = T522 ? 6'h28 : T493;
  assign T493 = T521 ? 6'h29 : T494;
  assign T494 = T520 ? 6'h2a : T495;
  assign T495 = T519 ? 6'h2b : T496;
  assign T496 = T518 ? 6'h2c : T497;
  assign T497 = T517 ? 6'h2d : T498;
  assign T498 = T516 ? 6'h2e : T499;
  assign T499 = T515 ? 6'h2f : T500;
  assign T500 = T514 ? 6'h30 : T501;
  assign T501 = T513 ? 6'h31 : T502;
  assign T502 = T503 ? 6'h32 : 6'h33;
  assign T503 = T12[50];
  assign T12 = {T50, T13};
  assign T13 = {T25, T14};
  assign T14 = {T21, T15};
  assign T15 = {T20, T16};
  assign T16 = T17[1];
  assign T17 = T18[3:2];
  assign T18 = T19[19:16];
  assign T19 = T7[51:32];
  assign T20 = T17[0];
  assign T21 = {T24, T22};
  assign T22 = T23[1];
  assign T23 = T18[1:0];
  assign T24 = T23[0];
  assign T25 = T48 | T26;
  assign T26 = T27 & 16'haaaa;
  assign T27 = T28 << 1'h1;
  assign T28 = T29[14:0];
  assign T29 = T46 | T30;
  assign T30 = T31 & 16'hcccc;
  assign T31 = T32 << 2'h2;
  assign T32 = T33[13:0];
  assign T33 = T44 | T34;
  assign T34 = T35 & 16'hf0f0;
  assign T35 = T36 << 3'h4;
  assign T36 = T37[11:0];
  assign T37 = T42 | T38;
  assign T38 = T39 & 16'hff00;
  assign T39 = T40 << 4'h8;
  assign T40 = T41[7:0];
  assign T41 = T19[15:0];
  assign T42 = T504 & 16'hff;
  assign T504 = {8'h0, T43};
  assign T43 = T41 >> 4'h8;
  assign T44 = T505 & 16'hf0f;
  assign T505 = {4'h0, T45};
  assign T45 = T37 >> 3'h4;
  assign T46 = T506 & 16'h3333;
  assign T506 = {2'h0, T47};
  assign T47 = T33 >> 2'h2;
  assign T48 = T507 & 16'h5555;
  assign T507 = {1'h0, T49};
  assign T49 = T29 >> 1'h1;
  assign T50 = T79 | T51;
  assign T51 = T52 & 32'haaaaaaaa;
  assign T52 = T53 << 1'h1;
  assign T53 = T54[30:0];
  assign T54 = T77 | T55;
  assign T55 = T56 & 32'hcccccccc;
  assign T56 = T57 << 2'h2;
  assign T57 = T58[29:0];
  assign T58 = T75 | T59;
  assign T59 = T60 & 32'hf0f0f0f0;
  assign T60 = T61 << 3'h4;
  assign T61 = T62[27:0];
  assign T62 = T73 | T63;
  assign T63 = T64 & 32'hff00ff00;
  assign T64 = T65 << 4'h8;
  assign T65 = T66[23:0];
  assign T66 = T71 | T67;
  assign T67 = T68 & 32'hffff0000;
  assign T68 = T69 << 5'h10;
  assign T69 = T70[15:0];
  assign T70 = T7[31:0];
  assign T71 = T508 & 32'hffff;
  assign T508 = {16'h0, T72};
  assign T72 = T70 >> 5'h10;
  assign T73 = T509 & 32'hff00ff;
  assign T509 = {8'h0, T74};
  assign T74 = T66 >> 4'h8;
  assign T75 = T510 & 32'hf0f0f0f;
  assign T510 = {4'h0, T76};
  assign T76 = T62 >> 3'h4;
  assign T77 = T511 & 32'h33333333;
  assign T511 = {2'h0, T78};
  assign T78 = T58 >> 2'h2;
  assign T79 = T512 & 32'h55555555;
  assign T512 = {1'h0, T80};
  assign T80 = T54 >> 1'h1;
  assign T513 = T12[49];
  assign T514 = T12[48];
  assign T515 = T12[47];
  assign T516 = T12[46];
  assign T517 = T12[45];
  assign T518 = T12[44];
  assign T519 = T12[43];
  assign T520 = T12[42];
  assign T521 = T12[41];
  assign T522 = T12[40];
  assign T523 = T12[39];
  assign T524 = T12[38];
  assign T525 = T12[37];
  assign T526 = T12[36];
  assign T527 = T12[35];
  assign T528 = T12[34];
  assign T529 = T12[33];
  assign T530 = T12[32];
  assign T531 = T12[31];
  assign T532 = T12[30];
  assign T533 = T12[29];
  assign T534 = T12[28];
  assign T535 = T12[27];
  assign T536 = T12[26];
  assign T537 = T12[25];
  assign T538 = T12[24];
  assign T539 = T12[23];
  assign T540 = T12[22];
  assign T541 = T12[21];
  assign T542 = T12[20];
  assign T543 = T12[19];
  assign T544 = T12[18];
  assign T545 = T12[17];
  assign T546 = T12[16];
  assign T547 = T12[15];
  assign T548 = T12[14];
  assign T549 = T12[13];
  assign T550 = T12[12];
  assign T551 = T12[11];
  assign T552 = T12[10];
  assign T553 = T12[9];
  assign T554 = T12[8];
  assign T555 = T12[7];
  assign T556 = T12[6];
  assign T557 = T12[5];
  assign T558 = T12[4];
  assign T559 = T12[3];
  assign T560 = T12[2];
  assign T561 = T12[1];
  assign T562 = T12[0];
  assign T81 = T82 == 11'h0;
  assign T82 = io_c[62:52];
  assign T83 = T84 ^ 1'h1;
  assign T84 = T81 & T85;
  assign T85 = T7 == 52'h0;
  assign T86 = T87[8:0];
  assign T87 = T88;
  assign T88 = T89;
  assign T89 = {1'h0, T90};
  assign T90 = T91;
  assign T91 = T94 + T563;
  assign T563 = {1'h0, T92};
  assign T92 = 11'h400 | T564;
  assign T564 = {9'h0, T93};
  assign T93 = T81 ? 2'h2 : 2'h1;
  assign T94 = T81 ? T95 : T565;
  assign T565 = {1'h0, T82};
  assign T95 = T566 ^ 12'hfff;
  assign T566 = {6'h0, T452};
  assign T96 = {T106, T97};
  assign T97 = T103 | T567;
  assign T567 = {2'h0, T98};
  assign T98 = T99;
  assign T99 = T101 & T100;
  assign T100 = T85 ^ 1'h1;
  assign T101 = T102 == 2'h3;
  assign T102 = T91[11:10];
  assign T103 = T105 ? 3'h0 : T104;
  assign T104 = T87[11:9];
  assign T105 = T84;
  assign T106 = T107;
  assign T107 = io_c[63];
  assign T108 = {T204, T109};
  assign T109 = {T194, T110};
  assign T110 = T111[51:0];
  assign T111 = T112;
  assign T112 = {1'h0, T113};
  assign T113 = {T191, T114};
  assign T114 = T189 ? T116 : T115;
  assign T115 = io_b[51:0];
  assign T116 = T117 << 1'h1;
  assign T117 = T118[50:0];
  assign T118 = T115 << T568;
  assign T568 = T678 ? 1'h0 : T569;
  assign T569 = T677 ? 1'h1 : T570;
  assign T570 = T676 ? 2'h2 : T571;
  assign T571 = T675 ? 2'h3 : T572;
  assign T572 = T674 ? 3'h4 : T573;
  assign T573 = T673 ? 3'h5 : T574;
  assign T574 = T672 ? 3'h6 : T575;
  assign T575 = T671 ? 3'h7 : T576;
  assign T576 = T670 ? 4'h8 : T577;
  assign T577 = T669 ? 4'h9 : T578;
  assign T578 = T668 ? 4'ha : T579;
  assign T579 = T667 ? 4'hb : T580;
  assign T580 = T666 ? 4'hc : T581;
  assign T581 = T665 ? 4'hd : T582;
  assign T582 = T664 ? 4'he : T583;
  assign T583 = T663 ? 4'hf : T584;
  assign T584 = T662 ? 5'h10 : T585;
  assign T585 = T661 ? 5'h11 : T586;
  assign T586 = T660 ? 5'h12 : T587;
  assign T587 = T659 ? 5'h13 : T588;
  assign T588 = T658 ? 5'h14 : T589;
  assign T589 = T657 ? 5'h15 : T590;
  assign T590 = T656 ? 5'h16 : T591;
  assign T591 = T655 ? 5'h17 : T592;
  assign T592 = T654 ? 5'h18 : T593;
  assign T593 = T653 ? 5'h19 : T594;
  assign T594 = T652 ? 5'h1a : T595;
  assign T595 = T651 ? 5'h1b : T596;
  assign T596 = T650 ? 5'h1c : T597;
  assign T597 = T649 ? 5'h1d : T598;
  assign T598 = T648 ? 5'h1e : T599;
  assign T599 = T647 ? 5'h1f : T600;
  assign T600 = T646 ? 6'h20 : T601;
  assign T601 = T645 ? 6'h21 : T602;
  assign T602 = T644 ? 6'h22 : T603;
  assign T603 = T643 ? 6'h23 : T604;
  assign T604 = T642 ? 6'h24 : T605;
  assign T605 = T641 ? 6'h25 : T606;
  assign T606 = T640 ? 6'h26 : T607;
  assign T607 = T639 ? 6'h27 : T608;
  assign T608 = T638 ? 6'h28 : T609;
  assign T609 = T637 ? 6'h29 : T610;
  assign T610 = T636 ? 6'h2a : T611;
  assign T611 = T635 ? 6'h2b : T612;
  assign T612 = T634 ? 6'h2c : T613;
  assign T613 = T633 ? 6'h2d : T614;
  assign T614 = T632 ? 6'h2e : T615;
  assign T615 = T631 ? 6'h2f : T616;
  assign T616 = T630 ? 6'h30 : T617;
  assign T617 = T629 ? 6'h31 : T618;
  assign T618 = T619 ? 6'h32 : 6'h33;
  assign T619 = T120[50];
  assign T120 = {T158, T121};
  assign T121 = {T133, T122};
  assign T122 = {T129, T123};
  assign T123 = {T128, T124};
  assign T124 = T125[1];
  assign T125 = T126[3:2];
  assign T126 = T127[19:16];
  assign T127 = T115[51:32];
  assign T128 = T125[0];
  assign T129 = {T132, T130};
  assign T130 = T131[1];
  assign T131 = T126[1:0];
  assign T132 = T131[0];
  assign T133 = T156 | T134;
  assign T134 = T135 & 16'haaaa;
  assign T135 = T136 << 1'h1;
  assign T136 = T137[14:0];
  assign T137 = T154 | T138;
  assign T138 = T139 & 16'hcccc;
  assign T139 = T140 << 2'h2;
  assign T140 = T141[13:0];
  assign T141 = T152 | T142;
  assign T142 = T143 & 16'hf0f0;
  assign T143 = T144 << 3'h4;
  assign T144 = T145[11:0];
  assign T145 = T150 | T146;
  assign T146 = T147 & 16'hff00;
  assign T147 = T148 << 4'h8;
  assign T148 = T149[7:0];
  assign T149 = T127[15:0];
  assign T150 = T620 & 16'hff;
  assign T620 = {8'h0, T151};
  assign T151 = T149 >> 4'h8;
  assign T152 = T621 & 16'hf0f;
  assign T621 = {4'h0, T153};
  assign T153 = T145 >> 3'h4;
  assign T154 = T622 & 16'h3333;
  assign T622 = {2'h0, T155};
  assign T155 = T141 >> 2'h2;
  assign T156 = T623 & 16'h5555;
  assign T623 = {1'h0, T157};
  assign T157 = T137 >> 1'h1;
  assign T158 = T187 | T159;
  assign T159 = T160 & 32'haaaaaaaa;
  assign T160 = T161 << 1'h1;
  assign T161 = T162[30:0];
  assign T162 = T185 | T163;
  assign T163 = T164 & 32'hcccccccc;
  assign T164 = T165 << 2'h2;
  assign T165 = T166[29:0];
  assign T166 = T183 | T167;
  assign T167 = T168 & 32'hf0f0f0f0;
  assign T168 = T169 << 3'h4;
  assign T169 = T170[27:0];
  assign T170 = T181 | T171;
  assign T171 = T172 & 32'hff00ff00;
  assign T172 = T173 << 4'h8;
  assign T173 = T174[23:0];
  assign T174 = T179 | T175;
  assign T175 = T176 & 32'hffff0000;
  assign T176 = T177 << 5'h10;
  assign T177 = T178[15:0];
  assign T178 = T115[31:0];
  assign T179 = T624 & 32'hffff;
  assign T624 = {16'h0, T180};
  assign T180 = T178 >> 5'h10;
  assign T181 = T625 & 32'hff00ff;
  assign T625 = {8'h0, T182};
  assign T182 = T174 >> 4'h8;
  assign T183 = T626 & 32'hf0f0f0f;
  assign T626 = {4'h0, T184};
  assign T184 = T170 >> 3'h4;
  assign T185 = T627 & 32'h33333333;
  assign T627 = {2'h0, T186};
  assign T186 = T166 >> 2'h2;
  assign T187 = T628 & 32'h55555555;
  assign T628 = {1'h0, T188};
  assign T188 = T162 >> 1'h1;
  assign T629 = T120[49];
  assign T630 = T120[48];
  assign T631 = T120[47];
  assign T632 = T120[46];
  assign T633 = T120[45];
  assign T634 = T120[44];
  assign T635 = T120[43];
  assign T636 = T120[42];
  assign T637 = T120[41];
  assign T638 = T120[40];
  assign T639 = T120[39];
  assign T640 = T120[38];
  assign T641 = T120[37];
  assign T642 = T120[36];
  assign T643 = T120[35];
  assign T644 = T120[34];
  assign T645 = T120[33];
  assign T646 = T120[32];
  assign T647 = T120[31];
  assign T648 = T120[30];
  assign T649 = T120[29];
  assign T650 = T120[28];
  assign T651 = T120[27];
  assign T652 = T120[26];
  assign T653 = T120[25];
  assign T654 = T120[24];
  assign T655 = T120[23];
  assign T656 = T120[22];
  assign T657 = T120[21];
  assign T658 = T120[20];
  assign T659 = T120[19];
  assign T660 = T120[18];
  assign T661 = T120[17];
  assign T662 = T120[16];
  assign T663 = T120[15];
  assign T664 = T120[14];
  assign T665 = T120[13];
  assign T666 = T120[12];
  assign T667 = T120[11];
  assign T668 = T120[10];
  assign T669 = T120[9];
  assign T670 = T120[8];
  assign T671 = T120[7];
  assign T672 = T120[6];
  assign T673 = T120[5];
  assign T674 = T120[4];
  assign T675 = T120[3];
  assign T676 = T120[2];
  assign T677 = T120[1];
  assign T678 = T120[0];
  assign T189 = T190 == 11'h0;
  assign T190 = io_b[62:52];
  assign T191 = T192 ^ 1'h1;
  assign T192 = T189 & T193;
  assign T193 = T115 == 52'h0;
  assign T194 = T195[8:0];
  assign T195 = T196;
  assign T196 = T197;
  assign T197 = {1'h0, T198};
  assign T198 = T199;
  assign T199 = T202 + T679;
  assign T679 = {1'h0, T200};
  assign T200 = 11'h400 | T680;
  assign T680 = {9'h0, T201};
  assign T201 = T189 ? 2'h2 : 2'h1;
  assign T202 = T189 ? T203 : T681;
  assign T681 = {1'h0, T190};
  assign T203 = T682 ^ 12'hfff;
  assign T682 = {6'h0, T568};
  assign T204 = {T214, T205};
  assign T205 = T211 | T683;
  assign T683 = {2'h0, T206};
  assign T206 = T207;
  assign T207 = T209 & T208;
  assign T208 = T193 ^ 1'h1;
  assign T209 = T210 == 2'h3;
  assign T210 = T199[11:10];
  assign T211 = T213 ? 3'h0 : T212;
  assign T212 = T195[11:9];
  assign T213 = T192;
  assign T214 = T215;
  assign T215 = io_b[63];
  assign T216 = {T312, T217};
  assign T217 = {T302, T218};
  assign T218 = T219[51:0];
  assign T219 = T220;
  assign T220 = {1'h0, T221};
  assign T221 = {T299, T222};
  assign T222 = T297 ? T224 : T223;
  assign T223 = io_a[51:0];
  assign T224 = T225 << 1'h1;
  assign T225 = T226[50:0];
  assign T226 = T223 << T684;
  assign T684 = T794 ? 1'h0 : T685;
  assign T685 = T793 ? 1'h1 : T686;
  assign T686 = T792 ? 2'h2 : T687;
  assign T687 = T791 ? 2'h3 : T688;
  assign T688 = T790 ? 3'h4 : T689;
  assign T689 = T789 ? 3'h5 : T690;
  assign T690 = T788 ? 3'h6 : T691;
  assign T691 = T787 ? 3'h7 : T692;
  assign T692 = T786 ? 4'h8 : T693;
  assign T693 = T785 ? 4'h9 : T694;
  assign T694 = T784 ? 4'ha : T695;
  assign T695 = T783 ? 4'hb : T696;
  assign T696 = T782 ? 4'hc : T697;
  assign T697 = T781 ? 4'hd : T698;
  assign T698 = T780 ? 4'he : T699;
  assign T699 = T779 ? 4'hf : T700;
  assign T700 = T778 ? 5'h10 : T701;
  assign T701 = T777 ? 5'h11 : T702;
  assign T702 = T776 ? 5'h12 : T703;
  assign T703 = T775 ? 5'h13 : T704;
  assign T704 = T774 ? 5'h14 : T705;
  assign T705 = T773 ? 5'h15 : T706;
  assign T706 = T772 ? 5'h16 : T707;
  assign T707 = T771 ? 5'h17 : T708;
  assign T708 = T770 ? 5'h18 : T709;
  assign T709 = T769 ? 5'h19 : T710;
  assign T710 = T768 ? 5'h1a : T711;
  assign T711 = T767 ? 5'h1b : T712;
  assign T712 = T766 ? 5'h1c : T713;
  assign T713 = T765 ? 5'h1d : T714;
  assign T714 = T764 ? 5'h1e : T715;
  assign T715 = T763 ? 5'h1f : T716;
  assign T716 = T762 ? 6'h20 : T717;
  assign T717 = T761 ? 6'h21 : T718;
  assign T718 = T760 ? 6'h22 : T719;
  assign T719 = T759 ? 6'h23 : T720;
  assign T720 = T758 ? 6'h24 : T721;
  assign T721 = T757 ? 6'h25 : T722;
  assign T722 = T756 ? 6'h26 : T723;
  assign T723 = T755 ? 6'h27 : T724;
  assign T724 = T754 ? 6'h28 : T725;
  assign T725 = T753 ? 6'h29 : T726;
  assign T726 = T752 ? 6'h2a : T727;
  assign T727 = T751 ? 6'h2b : T728;
  assign T728 = T750 ? 6'h2c : T729;
  assign T729 = T749 ? 6'h2d : T730;
  assign T730 = T748 ? 6'h2e : T731;
  assign T731 = T747 ? 6'h2f : T732;
  assign T732 = T746 ? 6'h30 : T733;
  assign T733 = T745 ? 6'h31 : T734;
  assign T734 = T735 ? 6'h32 : 6'h33;
  assign T735 = T228[50];
  assign T228 = {T266, T229};
  assign T229 = {T241, T230};
  assign T230 = {T237, T231};
  assign T231 = {T236, T232};
  assign T232 = T233[1];
  assign T233 = T234[3:2];
  assign T234 = T235[19:16];
  assign T235 = T223[51:32];
  assign T236 = T233[0];
  assign T237 = {T240, T238};
  assign T238 = T239[1];
  assign T239 = T234[1:0];
  assign T240 = T239[0];
  assign T241 = T264 | T242;
  assign T242 = T243 & 16'haaaa;
  assign T243 = T244 << 1'h1;
  assign T244 = T245[14:0];
  assign T245 = T262 | T246;
  assign T246 = T247 & 16'hcccc;
  assign T247 = T248 << 2'h2;
  assign T248 = T249[13:0];
  assign T249 = T260 | T250;
  assign T250 = T251 & 16'hf0f0;
  assign T251 = T252 << 3'h4;
  assign T252 = T253[11:0];
  assign T253 = T258 | T254;
  assign T254 = T255 & 16'hff00;
  assign T255 = T256 << 4'h8;
  assign T256 = T257[7:0];
  assign T257 = T235[15:0];
  assign T258 = T736 & 16'hff;
  assign T736 = {8'h0, T259};
  assign T259 = T257 >> 4'h8;
  assign T260 = T737 & 16'hf0f;
  assign T737 = {4'h0, T261};
  assign T261 = T253 >> 3'h4;
  assign T262 = T738 & 16'h3333;
  assign T738 = {2'h0, T263};
  assign T263 = T249 >> 2'h2;
  assign T264 = T739 & 16'h5555;
  assign T739 = {1'h0, T265};
  assign T265 = T245 >> 1'h1;
  assign T266 = T295 | T267;
  assign T267 = T268 & 32'haaaaaaaa;
  assign T268 = T269 << 1'h1;
  assign T269 = T270[30:0];
  assign T270 = T293 | T271;
  assign T271 = T272 & 32'hcccccccc;
  assign T272 = T273 << 2'h2;
  assign T273 = T274[29:0];
  assign T274 = T291 | T275;
  assign T275 = T276 & 32'hf0f0f0f0;
  assign T276 = T277 << 3'h4;
  assign T277 = T278[27:0];
  assign T278 = T289 | T279;
  assign T279 = T280 & 32'hff00ff00;
  assign T280 = T281 << 4'h8;
  assign T281 = T282[23:0];
  assign T282 = T287 | T283;
  assign T283 = T284 & 32'hffff0000;
  assign T284 = T285 << 5'h10;
  assign T285 = T286[15:0];
  assign T286 = T223[31:0];
  assign T287 = T740 & 32'hffff;
  assign T740 = {16'h0, T288};
  assign T288 = T286 >> 5'h10;
  assign T289 = T741 & 32'hff00ff;
  assign T741 = {8'h0, T290};
  assign T290 = T282 >> 4'h8;
  assign T291 = T742 & 32'hf0f0f0f;
  assign T742 = {4'h0, T292};
  assign T292 = T278 >> 3'h4;
  assign T293 = T743 & 32'h33333333;
  assign T743 = {2'h0, T294};
  assign T294 = T274 >> 2'h2;
  assign T295 = T744 & 32'h55555555;
  assign T744 = {1'h0, T296};
  assign T296 = T270 >> 1'h1;
  assign T745 = T228[49];
  assign T746 = T228[48];
  assign T747 = T228[47];
  assign T748 = T228[46];
  assign T749 = T228[45];
  assign T750 = T228[44];
  assign T751 = T228[43];
  assign T752 = T228[42];
  assign T753 = T228[41];
  assign T754 = T228[40];
  assign T755 = T228[39];
  assign T756 = T228[38];
  assign T757 = T228[37];
  assign T758 = T228[36];
  assign T759 = T228[35];
  assign T760 = T228[34];
  assign T761 = T228[33];
  assign T762 = T228[32];
  assign T763 = T228[31];
  assign T764 = T228[30];
  assign T765 = T228[29];
  assign T766 = T228[28];
  assign T767 = T228[27];
  assign T768 = T228[26];
  assign T769 = T228[25];
  assign T770 = T228[24];
  assign T771 = T228[23];
  assign T772 = T228[22];
  assign T773 = T228[21];
  assign T774 = T228[20];
  assign T775 = T228[19];
  assign T776 = T228[18];
  assign T777 = T228[17];
  assign T778 = T228[16];
  assign T779 = T228[15];
  assign T780 = T228[14];
  assign T781 = T228[13];
  assign T782 = T228[12];
  assign T783 = T228[11];
  assign T784 = T228[10];
  assign T785 = T228[9];
  assign T786 = T228[8];
  assign T787 = T228[7];
  assign T788 = T228[6];
  assign T789 = T228[5];
  assign T790 = T228[4];
  assign T791 = T228[3];
  assign T792 = T228[2];
  assign T793 = T228[1];
  assign T794 = T228[0];
  assign T297 = T298 == 11'h0;
  assign T298 = io_a[62:52];
  assign T299 = T300 ^ 1'h1;
  assign T300 = T297 & T301;
  assign T301 = T223 == 52'h0;
  assign T302 = T303[8:0];
  assign T303 = T304;
  assign T304 = T305;
  assign T305 = {1'h0, T306};
  assign T306 = T307;
  assign T307 = T310 + T795;
  assign T795 = {1'h0, T308};
  assign T308 = 11'h400 | T796;
  assign T796 = {9'h0, T309};
  assign T309 = T297 ? 2'h2 : 2'h1;
  assign T310 = T297 ? T311 : T797;
  assign T797 = {1'h0, T298};
  assign T311 = T798 ^ 12'hfff;
  assign T798 = {6'h0, T684};
  assign T312 = {T322, T313};
  assign T313 = T319 | T799;
  assign T799 = {2'h0, T314};
  assign T314 = T315;
  assign T315 = T317 & T316;
  assign T316 = T301 ^ 1'h1;
  assign T317 = T318 == 2'h3;
  assign T318 = T307[11:10];
  assign T319 = T321 ? 3'h0 : T320;
  assign T320 = T303[11:9];
  assign T321 = T300;
  assign T322 = T323;
  assign T323 = io_a[63];
  assign io_pass = T324;
  assign T324 = T326 & T325;
  assign T325 = io_actual_exceptionFlags == io_expected_exceptionFlags;
  assign T326 = T339 ? T334 : T327;
  assign T327 = T332 ? T329 : T328;
  assign T328 = io_actual_out == io_expected_recOut;
  assign T329 = T331 == T330;
  assign T330 = io_expected_recOut[64:61];
  assign T331 = io_actual_out[64:61];
  assign T332 = T333 == 3'h6;
  assign T333 = T331[2:0];
  assign T334 = T338 & T335;
  assign T335 = T337 == T336;
  assign T336 = io_expected_recOut[51:0];
  assign T337 = io_actual_out[51:0];
  assign T338 = T331 == T330;
  assign T339 = T342 | T340;
  assign T340 = T341 == 3'h7;
  assign T341 = T331[2:0];
  assign T342 = T343 == 3'h0;
  assign T343 = T331[2:0];
  assign io_check = 1'h1;
  assign io_actual_exceptionFlags = mulAddRecFN_io_exceptionFlags;
  assign io_actual_out = mulAddRecFN_io_out;
  assign io_expected_recOut = T344;
  assign T344 = {T440, T345};
  assign T345 = {T430, T346};
  assign T346 = T347[51:0];
  assign T347 = T348;
  assign T348 = {1'h0, T349};
  assign T349 = {T427, T350};
  assign T350 = T425 ? T352 : T351;
  assign T351 = io_expected_out[51:0];
  assign T352 = T353 << 1'h1;
  assign T353 = T354[50:0];
  assign T354 = T351 << T800;
  assign T800 = T910 ? 1'h0 : T801;
  assign T801 = T909 ? 1'h1 : T802;
  assign T802 = T908 ? 2'h2 : T803;
  assign T803 = T907 ? 2'h3 : T804;
  assign T804 = T906 ? 3'h4 : T805;
  assign T805 = T905 ? 3'h5 : T806;
  assign T806 = T904 ? 3'h6 : T807;
  assign T807 = T903 ? 3'h7 : T808;
  assign T808 = T902 ? 4'h8 : T809;
  assign T809 = T901 ? 4'h9 : T810;
  assign T810 = T900 ? 4'ha : T811;
  assign T811 = T899 ? 4'hb : T812;
  assign T812 = T898 ? 4'hc : T813;
  assign T813 = T897 ? 4'hd : T814;
  assign T814 = T896 ? 4'he : T815;
  assign T815 = T895 ? 4'hf : T816;
  assign T816 = T894 ? 5'h10 : T817;
  assign T817 = T893 ? 5'h11 : T818;
  assign T818 = T892 ? 5'h12 : T819;
  assign T819 = T891 ? 5'h13 : T820;
  assign T820 = T890 ? 5'h14 : T821;
  assign T821 = T889 ? 5'h15 : T822;
  assign T822 = T888 ? 5'h16 : T823;
  assign T823 = T887 ? 5'h17 : T824;
  assign T824 = T886 ? 5'h18 : T825;
  assign T825 = T885 ? 5'h19 : T826;
  assign T826 = T884 ? 5'h1a : T827;
  assign T827 = T883 ? 5'h1b : T828;
  assign T828 = T882 ? 5'h1c : T829;
  assign T829 = T881 ? 5'h1d : T830;
  assign T830 = T880 ? 5'h1e : T831;
  assign T831 = T879 ? 5'h1f : T832;
  assign T832 = T878 ? 6'h20 : T833;
  assign T833 = T877 ? 6'h21 : T834;
  assign T834 = T876 ? 6'h22 : T835;
  assign T835 = T875 ? 6'h23 : T836;
  assign T836 = T874 ? 6'h24 : T837;
  assign T837 = T873 ? 6'h25 : T838;
  assign T838 = T872 ? 6'h26 : T839;
  assign T839 = T871 ? 6'h27 : T840;
  assign T840 = T870 ? 6'h28 : T841;
  assign T841 = T869 ? 6'h29 : T842;
  assign T842 = T868 ? 6'h2a : T843;
  assign T843 = T867 ? 6'h2b : T844;
  assign T844 = T866 ? 6'h2c : T845;
  assign T845 = T865 ? 6'h2d : T846;
  assign T846 = T864 ? 6'h2e : T847;
  assign T847 = T863 ? 6'h2f : T848;
  assign T848 = T862 ? 6'h30 : T849;
  assign T849 = T861 ? 6'h31 : T850;
  assign T850 = T851 ? 6'h32 : 6'h33;
  assign T851 = T356[50];
  assign T356 = {T394, T357};
  assign T357 = {T369, T358};
  assign T358 = {T365, T359};
  assign T359 = {T364, T360};
  assign T360 = T361[1];
  assign T361 = T362[3:2];
  assign T362 = T363[19:16];
  assign T363 = T351[51:32];
  assign T364 = T361[0];
  assign T365 = {T368, T366};
  assign T366 = T367[1];
  assign T367 = T362[1:0];
  assign T368 = T367[0];
  assign T369 = T392 | T370;
  assign T370 = T371 & 16'haaaa;
  assign T371 = T372 << 1'h1;
  assign T372 = T373[14:0];
  assign T373 = T390 | T374;
  assign T374 = T375 & 16'hcccc;
  assign T375 = T376 << 2'h2;
  assign T376 = T377[13:0];
  assign T377 = T388 | T378;
  assign T378 = T379 & 16'hf0f0;
  assign T379 = T380 << 3'h4;
  assign T380 = T381[11:0];
  assign T381 = T386 | T382;
  assign T382 = T383 & 16'hff00;
  assign T383 = T384 << 4'h8;
  assign T384 = T385[7:0];
  assign T385 = T363[15:0];
  assign T386 = T852 & 16'hff;
  assign T852 = {8'h0, T387};
  assign T387 = T385 >> 4'h8;
  assign T388 = T853 & 16'hf0f;
  assign T853 = {4'h0, T389};
  assign T389 = T381 >> 3'h4;
  assign T390 = T854 & 16'h3333;
  assign T854 = {2'h0, T391};
  assign T391 = T377 >> 2'h2;
  assign T392 = T855 & 16'h5555;
  assign T855 = {1'h0, T393};
  assign T393 = T373 >> 1'h1;
  assign T394 = T423 | T395;
  assign T395 = T396 & 32'haaaaaaaa;
  assign T396 = T397 << 1'h1;
  assign T397 = T398[30:0];
  assign T398 = T421 | T399;
  assign T399 = T400 & 32'hcccccccc;
  assign T400 = T401 << 2'h2;
  assign T401 = T402[29:0];
  assign T402 = T419 | T403;
  assign T403 = T404 & 32'hf0f0f0f0;
  assign T404 = T405 << 3'h4;
  assign T405 = T406[27:0];
  assign T406 = T417 | T407;
  assign T407 = T408 & 32'hff00ff00;
  assign T408 = T409 << 4'h8;
  assign T409 = T410[23:0];
  assign T410 = T415 | T411;
  assign T411 = T412 & 32'hffff0000;
  assign T412 = T413 << 5'h10;
  assign T413 = T414[15:0];
  assign T414 = T351[31:0];
  assign T415 = T856 & 32'hffff;
  assign T856 = {16'h0, T416};
  assign T416 = T414 >> 5'h10;
  assign T417 = T857 & 32'hff00ff;
  assign T857 = {8'h0, T418};
  assign T418 = T410 >> 4'h8;
  assign T419 = T858 & 32'hf0f0f0f;
  assign T858 = {4'h0, T420};
  assign T420 = T406 >> 3'h4;
  assign T421 = T859 & 32'h33333333;
  assign T859 = {2'h0, T422};
  assign T422 = T402 >> 2'h2;
  assign T423 = T860 & 32'h55555555;
  assign T860 = {1'h0, T424};
  assign T424 = T398 >> 1'h1;
  assign T861 = T356[49];
  assign T862 = T356[48];
  assign T863 = T356[47];
  assign T864 = T356[46];
  assign T865 = T356[45];
  assign T866 = T356[44];
  assign T867 = T356[43];
  assign T868 = T356[42];
  assign T869 = T356[41];
  assign T870 = T356[40];
  assign T871 = T356[39];
  assign T872 = T356[38];
  assign T873 = T356[37];
  assign T874 = T356[36];
  assign T875 = T356[35];
  assign T876 = T356[34];
  assign T877 = T356[33];
  assign T878 = T356[32];
  assign T879 = T356[31];
  assign T880 = T356[30];
  assign T881 = T356[29];
  assign T882 = T356[28];
  assign T883 = T356[27];
  assign T884 = T356[26];
  assign T885 = T356[25];
  assign T886 = T356[24];
  assign T887 = T356[23];
  assign T888 = T356[22];
  assign T889 = T356[21];
  assign T890 = T356[20];
  assign T891 = T356[19];
  assign T892 = T356[18];
  assign T893 = T356[17];
  assign T894 = T356[16];
  assign T895 = T356[15];
  assign T896 = T356[14];
  assign T897 = T356[13];
  assign T898 = T356[12];
  assign T899 = T356[11];
  assign T900 = T356[10];
  assign T901 = T356[9];
  assign T902 = T356[8];
  assign T903 = T356[7];
  assign T904 = T356[6];
  assign T905 = T356[5];
  assign T906 = T356[4];
  assign T907 = T356[3];
  assign T908 = T356[2];
  assign T909 = T356[1];
  assign T910 = T356[0];
  assign T425 = T426 == 11'h0;
  assign T426 = io_expected_out[62:52];
  assign T427 = T428 ^ 1'h1;
  assign T428 = T425 & T429;
  assign T429 = T351 == 52'h0;
  assign T430 = T431[8:0];
  assign T431 = T432;
  assign T432 = T433;
  assign T433 = {1'h0, T434};
  assign T434 = T435;
  assign T435 = T438 + T911;
  assign T911 = {1'h0, T436};
  assign T436 = 11'h400 | T912;
  assign T912 = {9'h0, T437};
  assign T437 = T425 ? 2'h2 : 2'h1;
  assign T438 = T425 ? T439 : T913;
  assign T913 = {1'h0, T426};
  assign T439 = T914 ^ 12'hfff;
  assign T914 = {6'h0, T800};
  assign T440 = {T450, T441};
  assign T441 = T447 | T915;
  assign T915 = {2'h0, T442};
  assign T442 = T443;
  assign T443 = T445 & T444;
  assign T444 = T429 ^ 1'h1;
  assign T445 = T446 == 2'h3;
  assign T446 = T435[11:10];
  assign T447 = T449 ? 3'h0 : T448;
  assign T448 = T431[11:9];
  assign T449 = T428;
  assign T450 = T451;
  assign T451 = io_expected_out[63];
  MulAddRecFN mulAddRecFN(
       .io_op( 2'h0 ),
       .io_a( T216 ),
       .io_b( T108 ),
       .io_c( T0 ),
       .io_roundingMode( io_roundingMode ),
       .io_detectTininess( io_detectTininess ),
       .io_out( mulAddRecFN_io_out ),
       .io_exceptionFlags( mulAddRecFN_io_exceptionFlags )
  );
endmodule

