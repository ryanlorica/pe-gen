module MulAddRecFNToRaw_preMul(
    input [1:0] io_op,
    input [64:0] io_a,
    input [64:0] io_b,
    input [64:0] io_c,
    output[52:0] io_mulAddA,
    output[52:0] io_mulAddB,
    output[105:0] io_mulAddC,
    output io_toPostMul_isSigNaNAny,
    output io_toPostMul_isNaNAOrB,
    output io_toPostMul_isInfA,
    output io_toPostMul_isZeroA,
    output io_toPostMul_isInfB,
    output io_toPostMul_isZeroB,
    output io_toPostMul_signProd,
    output io_toPostMul_isNaNC,
    output io_toPostMul_isInfC,
    output io_toPostMul_isZeroC,
    output[12:0] io_toPostMul_sExpSum,
    output io_toPostMul_doSubMags,
    output io_toPostMul_CIsDominant,
    output[5:0] io_toPostMul_CDom_CAlignDist,
    output[54:0] io_toPostMul_highAlignedSigC,
    output io_toPostMul_bit0AlignedSigC
);

  wire T0;
  wire[162:0] alignedSigC;
  wire T1;
  wire T2;
  wire reduced4CExtra;
  wire[13:0] T3;
  wire[13:0] T190;
  wire[12:0] T4;
  wire[4:0] T5;
  wire T6;
  wire[4:0] T7;
  wire[12:0] T8;
  wire[64:0] T9;
  wire[5:0] T10;
  wire[7:0] CAlignDist;
  wire[7:0] T11;
  wire[7:0] T12;
  wire[12:0] posNatCAlignDist;
  wire[14:0] sNatCAlignDist;
  wire[13:0] T191;
  wire[12:0] rawC_sExp;
  wire[12:0] T13;
  wire[12:0] T14;
  wire[11:0] T15;
  wire T192;
  wire[14:0] sExpAlignedProd;
  wire[14:0] T16;
  wire[13:0] T193;
  wire[12:0] rawB_sExp;
  wire[12:0] T17;
  wire[12:0] T18;
  wire[11:0] T19;
  wire T194;
  wire[13:0] T195;
  wire[12:0] rawA_sExp;
  wire[12:0] T20;
  wire[12:0] T21;
  wire[11:0] T22;
  wire T196;
  wire T23;
  wire isMinCAlign;
  wire T24;
  wire T25;
  wire rawB_isZero;
  wire T26;
  wire[2:0] T27;
  wire rawA_isZero;
  wire T28;
  wire[2:0] T29;
  wire[3:0] T30;
  wire[1:0] T31;
  wire T32;
  wire[1:0] T33;
  wire[3:0] T34;
  wire T35;
  wire[1:0] T36;
  wire T37;
  wire[1:0] T38;
  wire T39;
  wire[7:0] T40;
  wire[7:0] T41;
  wire[7:0] T42;
  wire[6:0] T43;
  wire[7:0] T44;
  wire[7:0] T45;
  wire[7:0] T46;
  wire[5:0] T47;
  wire[7:0] T48;
  wire[7:0] T49;
  wire[7:0] T50;
  wire[3:0] T51;
  wire[7:0] T52;
  wire[7:0] T53;
  wire[7:0] T197;
  wire[3:0] T54;
  wire[7:0] T55;
  wire[7:0] T198;
  wire[5:0] T56;
  wire[7:0] T57;
  wire[7:0] T199;
  wire[6:0] T58;
  wire[13:0] T59;
  wire[13:0] T60;
  wire[6:0] T61;
  wire[3:0] T62;
  wire[1:0] T63;
  wire T64;
  wire T65;
  wire[3:0] T66;
  wire[53:0] T67;
  wire[53:0] rawC_sig;
  wire[53:0] T68;
  wire[52:0] T69;
  wire[51:0] T70;
  wire T71;
  wire T72;
  wire[2:0] T73;
  wire T74;
  wire T75;
  wire[3:0] T76;
  wire[1:0] T77;
  wire T78;
  wire T79;
  wire[3:0] T80;
  wire T81;
  wire T82;
  wire[3:0] T83;
  wire[2:0] T84;
  wire[1:0] T85;
  wire T86;
  wire T87;
  wire[3:0] T88;
  wire T89;
  wire T90;
  wire[3:0] T91;
  wire T92;
  wire T93;
  wire[3:0] T94;
  wire[6:0] T95;
  wire[3:0] T96;
  wire[1:0] T97;
  wire T98;
  wire T99;
  wire[3:0] T100;
  wire T101;
  wire T102;
  wire[3:0] T103;
  wire[1:0] T104;
  wire T105;
  wire T106;
  wire[3:0] T107;
  wire T108;
  wire T109;
  wire[3:0] T110;
  wire[2:0] T111;
  wire[1:0] T112;
  wire T113;
  wire T114;
  wire[3:0] T115;
  wire T116;
  wire T117;
  wire[3:0] T118;
  wire T119;
  wire T120;
  wire[1:0] T121;
  wire T122;
  wire[2:0] T123;
  wire[164:0] mainAlignedSigC;
  wire[164:0] T124;
  wire[164:0] T125;
  wire[110:0] T126;
  wire[110:0] T200;
  wire[53:0] T127;
  wire[53:0] T128;
  wire T129;
  wire T130;
  wire T131;
  wire[2:0] T132;
  wire doSubMags;
  wire T133;
  wire T134;
  wire rawC_sign;
  wire T135;
  wire signProd;
  wire T136;
  wire T137;
  wire rawB_sign;
  wire T138;
  wire rawA_sign;
  wire T139;
  wire[161:0] T140;
  wire[54:0] T141;
  wire[5:0] T142;
  wire CIsDominant;
  wire T143;
  wire T144;
  wire T145;
  wire rawC_isZero;
  wire[12:0] T201;
  wire[14:0] T146;
  wire[14:0] T147;
  wire[13:0] T202;
  wire T203;
  wire rawC_isInf;
  wire T148;
  wire T149;
  wire T150;
  wire T151;
  wire[1:0] T152;
  wire rawC_isNaN;
  wire T153;
  wire T154;
  wire rawB_isInf;
  wire T155;
  wire T156;
  wire T157;
  wire T158;
  wire[1:0] T159;
  wire rawA_isInf;
  wire T160;
  wire T161;
  wire T162;
  wire T163;
  wire[1:0] T164;
  wire T165;
  wire rawB_isNaN;
  wire T166;
  wire T167;
  wire rawA_isNaN;
  wire T168;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire T173;
  wire T174;
  wire T175;
  wire T176;
  wire T177;
  wire[53:0] rawB_sig;
  wire[53:0] T178;
  wire[52:0] T179;
  wire[51:0] T180;
  wire T181;
  wire T182;
  wire T183;
  wire T184;
  wire[53:0] rawA_sig;
  wire[53:0] T185;
  wire[52:0] T186;
  wire[51:0] T187;
  wire T188;
  wire[105:0] T189;
  wire[52:0] T204;
  wire[52:0] T205;


  assign io_toPostMul_bit0AlignedSigC = T0;
  assign T0 = alignedSigC[0];
  assign alignedSigC = {T140, T1};
  assign T1 = doSubMags ? T129 : T2;
  assign T2 = T122 | reduced4CExtra;
  assign reduced4CExtra = T3 != 14'h0;
  assign T3 = T59 & T190;
  assign T190 = {1'h0, T4};
  assign T4 = {T40, T5};
  assign T5 = {T30, T6};
  assign T6 = T7[4];
  assign T7 = T8[12:8];
  assign T8 = T9[36:24];
  assign T9 = $signed(65'h10000000000000000) >>> T10;
  assign T10 = CAlignDist >> 2'h2;
  assign CAlignDist = isMinCAlign ? 8'h0 : T11;
  assign T11 = T23 ? T12 : 8'ha1;
  assign T12 = posNatCAlignDist[7:0];
  assign posNatCAlignDist = sNatCAlignDist[12:0];
  assign sNatCAlignDist = sExpAlignedProd - T191;
  assign T191 = {T192, rawC_sExp};
  assign rawC_sExp = T13;
  assign T13 = T14;
  assign T14 = {1'h0, T15};
  assign T15 = io_c[63:52];
  assign T192 = rawC_sExp[12];
  assign sExpAlignedProd = T16 + 14'h3838;
  assign T16 = T195 + T193;
  assign T193 = {T194, rawB_sExp};
  assign rawB_sExp = T17;
  assign T17 = T18;
  assign T18 = {1'h0, T19};
  assign T19 = io_b[63:52];
  assign T194 = rawB_sExp[12];
  assign T195 = {T196, rawA_sExp};
  assign rawA_sExp = T20;
  assign T20 = T21;
  assign T21 = {1'h0, T22};
  assign T22 = io_a[63:52];
  assign T196 = rawA_sExp[12];
  assign T23 = posNatCAlignDist < 13'ha1;
  assign isMinCAlign = T25 | T24;
  assign T24 = $signed(sNatCAlignDist) < $signed(1'h0);
  assign T25 = rawA_isZero | rawB_isZero;
  assign rawB_isZero = T26;
  assign T26 = T27 == 3'h0;
  assign T27 = T19[11:9];
  assign rawA_isZero = T28;
  assign T28 = T29 == 3'h0;
  assign T29 = T22[11:9];
  assign T30 = {T36, T31};
  assign T31 = {T35, T32};
  assign T32 = T33[1];
  assign T33 = T34[3:2];
  assign T34 = T7[3:0];
  assign T35 = T33[0];
  assign T36 = {T39, T37};
  assign T37 = T38[1];
  assign T38 = T34[1:0];
  assign T39 = T38[0];
  assign T40 = T57 | T41;
  assign T41 = T42 & 8'haa;
  assign T42 = T43 << 1'h1;
  assign T43 = T44[6:0];
  assign T44 = T55 | T45;
  assign T45 = T46 & 8'hcc;
  assign T46 = T47 << 2'h2;
  assign T47 = T48[5:0];
  assign T48 = T53 | T49;
  assign T49 = T50 & 8'hf0;
  assign T50 = T51 << 3'h4;
  assign T51 = T52[3:0];
  assign T52 = T8[7:0];
  assign T53 = T197 & 8'hf;
  assign T197 = {4'h0, T54};
  assign T54 = T52 >> 3'h4;
  assign T55 = T198 & 8'h33;
  assign T198 = {2'h0, T56};
  assign T56 = T48 >> 2'h2;
  assign T57 = T199 & 8'h55;
  assign T199 = {1'h0, T58};
  assign T58 = T44 >> 1'h1;
  assign T59 = T60;
  assign T60 = {T95, T61};
  assign T61 = {T84, T62};
  assign T62 = {T77, T63};
  assign T63 = {T74, T64};
  assign T64 = T65;
  assign T65 = T66 != 4'h0;
  assign T66 = T67[3:0];
  assign T67 = rawC_sig << 1'h0;
  assign rawC_sig = T68;
  assign T68 = {1'h0, T69};
  assign T69 = {T71, T70};
  assign T70 = io_c[51:0];
  assign T71 = T72 ^ 1'h1;
  assign T72 = T73 == 3'h0;
  assign T73 = T15[11:9];
  assign T74 = T75;
  assign T75 = T76 != 4'h0;
  assign T76 = T67[7:4];
  assign T77 = {T81, T78};
  assign T78 = T79;
  assign T79 = T80 != 4'h0;
  assign T80 = T67[11:8];
  assign T81 = T82;
  assign T82 = T83 != 4'h0;
  assign T83 = T67[15:12];
  assign T84 = {T92, T85};
  assign T85 = {T89, T86};
  assign T86 = T87;
  assign T87 = T88 != 4'h0;
  assign T88 = T67[19:16];
  assign T89 = T90;
  assign T90 = T91 != 4'h0;
  assign T91 = T67[23:20];
  assign T92 = T93;
  assign T93 = T94 != 4'h0;
  assign T94 = T67[27:24];
  assign T95 = {T111, T96};
  assign T96 = {T104, T97};
  assign T97 = {T101, T98};
  assign T98 = T99;
  assign T99 = T100 != 4'h0;
  assign T100 = T67[31:28];
  assign T101 = T102;
  assign T102 = T103 != 4'h0;
  assign T103 = T67[35:32];
  assign T104 = {T108, T105};
  assign T105 = T106;
  assign T106 = T107 != 4'h0;
  assign T107 = T67[39:36];
  assign T108 = T109;
  assign T109 = T110 != 4'h0;
  assign T110 = T67[43:40];
  assign T111 = {T119, T112};
  assign T112 = {T116, T113};
  assign T113 = T114;
  assign T114 = T115 != 4'h0;
  assign T115 = T67[47:44];
  assign T116 = T117;
  assign T117 = T118 != 4'h0;
  assign T118 = T67[51:48];
  assign T119 = T120;
  assign T120 = T121 != 2'h0;
  assign T121 = T67[53:52];
  assign T122 = T123 != 3'h0;
  assign T123 = mainAlignedSigC[2:0];
  assign mainAlignedSigC = $signed(T124) >>> CAlignDist;
  assign T124 = T125;
  assign T125 = {T127, T126};
  assign T126 = 111'h0 - T200;
  assign T200 = {110'h0, doSubMags};
  assign T127 = doSubMags ? T128 : rawC_sig;
  assign T128 = ~ rawC_sig;
  assign T129 = T131 & T130;
  assign T130 = reduced4CExtra ^ 1'h1;
  assign T131 = T132 == 3'h7;
  assign T132 = mainAlignedSigC[2:0];
  assign doSubMags = T134 ^ T133;
  assign T133 = io_op[0];
  assign T134 = signProd ^ rawC_sign;
  assign rawC_sign = T135;
  assign T135 = io_c[64];
  assign signProd = T137 ^ T136;
  assign T136 = io_op[1];
  assign T137 = rawA_sign ^ rawB_sign;
  assign rawB_sign = T138;
  assign T138 = io_b[64];
  assign rawA_sign = T139;
  assign T139 = io_a[64];
  assign T140 = $signed(mainAlignedSigC) >>> 2'h3;
  assign io_toPostMul_highAlignedSigC = T141;
  assign T141 = alignedSigC[161:107];
  assign io_toPostMul_CDom_CAlignDist = T142;
  assign T142 = CAlignDist[5:0];
  assign io_toPostMul_CIsDominant = CIsDominant;
  assign CIsDominant = T145 & T143;
  assign T143 = isMinCAlign | T144;
  assign T144 = posNatCAlignDist <= 13'h35;
  assign T145 = rawC_isZero ^ 1'h1;
  assign rawC_isZero = T72;
  assign io_toPostMul_doSubMags = doSubMags;
  assign io_toPostMul_sExpSum = T201;
  assign T201 = T146[12:0];
  assign T146 = CIsDominant ? T202 : T147;
  assign T147 = sExpAlignedProd - 14'h35;
  assign T202 = {T203, rawC_sExp};
  assign T203 = rawC_sExp[12];
  assign io_toPostMul_isZeroC = rawC_isZero;
  assign io_toPostMul_isInfC = rawC_isInf;
  assign rawC_isInf = T148;
  assign T148 = T151 & T149;
  assign T149 = T150 ^ 1'h1;
  assign T150 = T15[9];
  assign T151 = T152 == 2'h3;
  assign T152 = T15[11:10];
  assign io_toPostMul_isNaNC = rawC_isNaN;
  assign rawC_isNaN = T153;
  assign T153 = T151 & T154;
  assign T154 = T15[9];
  assign io_toPostMul_signProd = signProd;
  assign io_toPostMul_isZeroB = rawB_isZero;
  assign io_toPostMul_isInfB = rawB_isInf;
  assign rawB_isInf = T155;
  assign T155 = T158 & T156;
  assign T156 = T157 ^ 1'h1;
  assign T157 = T19[9];
  assign T158 = T159 == 2'h3;
  assign T159 = T19[11:10];
  assign io_toPostMul_isZeroA = rawA_isZero;
  assign io_toPostMul_isInfA = rawA_isInf;
  assign rawA_isInf = T160;
  assign T160 = T163 & T161;
  assign T161 = T162 ^ 1'h1;
  assign T162 = T22[9];
  assign T163 = T164 == 2'h3;
  assign T164 = T22[11:10];
  assign io_toPostMul_isNaNAOrB = T165;
  assign T165 = rawA_isNaN | rawB_isNaN;
  assign rawB_isNaN = T166;
  assign T166 = T158 & T167;
  assign T167 = T19[9];
  assign rawA_isNaN = T168;
  assign T168 = T163 & T169;
  assign T169 = T22[9];
  assign io_toPostMul_isSigNaNAny = T170;
  assign T170 = T174 | T171;
  assign T171 = rawC_isNaN & T172;
  assign T172 = T173 ^ 1'h1;
  assign T173 = rawC_sig[51];
  assign T174 = T182 | T175;
  assign T175 = rawB_isNaN & T176;
  assign T176 = T177 ^ 1'h1;
  assign T177 = rawB_sig[51];
  assign rawB_sig = T178;
  assign T178 = {1'h0, T179};
  assign T179 = {T181, T180};
  assign T180 = io_b[51:0];
  assign T181 = T26 ^ 1'h1;
  assign T182 = rawA_isNaN & T183;
  assign T183 = T184 ^ 1'h1;
  assign T184 = rawA_sig[51];
  assign rawA_sig = T185;
  assign T185 = {1'h0, T186};
  assign T186 = {T188, T187};
  assign T187 = io_a[51:0];
  assign T188 = T28 ^ 1'h1;
  assign io_mulAddC = T189;
  assign T189 = alignedSigC[106:1];
  assign io_mulAddB = T204;
  assign T204 = rawB_sig[52:0];
  assign io_mulAddA = T205;
  assign T205 = rawA_sig[52:0];
endmodule

module MulAddRecFNToRaw_postMul(
    input  io_fromPreMul_isSigNaNAny,
    input  io_fromPreMul_isNaNAOrB,
    input  io_fromPreMul_isInfA,
    input  io_fromPreMul_isZeroA,
    input  io_fromPreMul_isInfB,
    input  io_fromPreMul_isZeroB,
    input  io_fromPreMul_signProd,
    input  io_fromPreMul_isNaNC,
    input  io_fromPreMul_isInfC,
    input  io_fromPreMul_isZeroC,
    input [12:0] io_fromPreMul_sExpSum,
    input  io_fromPreMul_doSubMags,
    input  io_fromPreMul_CIsDominant,
    input [5:0] io_fromPreMul_CDom_CAlignDist,
    input [54:0] io_fromPreMul_highAlignedSigC,
    input  io_fromPreMul_bit0AlignedSigC,
    input [106:0] io_mulAddResult,
    input [2:0] io_roundingMode,
    output io_invalidExc,
    output io_rawOut_isNaN,
    output io_rawOut_isInf,
    output io_rawOut_isZero,
    output io_rawOut_sign,
    output[12:0] io_rawOut_sExp,
    output[55:0] io_rawOut_sig
);

  wire[55:0] T0;
  wire[55:0] notCDom_sig;
  wire T1;
  wire notCDom_reduced4SigExtra;
  wire[13:0] T2;
  wire[13:0] T561;
  wire[12:0] T3;
  wire[4:0] T4;
  wire T5;
  wire[4:0] T6;
  wire[12:0] T7;
  wire[32:0] T8;
  wire[4:0] T9;
  wire[4:0] T10;
  wire[5:0] T562;
  wire[5:0] T563;
  wire[5:0] T564;
  wire[5:0] T565;
  wire[5:0] T566;
  wire[5:0] T567;
  wire[5:0] T568;
  wire[5:0] T569;
  wire[5:0] T570;
  wire[5:0] T571;
  wire[5:0] T572;
  wire[5:0] T573;
  wire[5:0] T574;
  wire[5:0] T575;
  wire[5:0] T576;
  wire[5:0] T577;
  wire[5:0] T578;
  wire[5:0] T579;
  wire[5:0] T580;
  wire[5:0] T581;
  wire[5:0] T582;
  wire[5:0] T583;
  wire[5:0] T584;
  wire[5:0] T585;
  wire[5:0] T586;
  wire[5:0] T587;
  wire[5:0] T588;
  wire[5:0] T589;
  wire[5:0] T590;
  wire[5:0] T591;
  wire[5:0] T592;
  wire[5:0] T593;
  wire[5:0] T594;
  wire[5:0] T595;
  wire[5:0] T596;
  wire[5:0] T597;
  wire[5:0] T598;
  wire[5:0] T599;
  wire[5:0] T600;
  wire[5:0] T601;
  wire[5:0] T602;
  wire[5:0] T603;
  wire[5:0] T604;
  wire[5:0] T605;
  wire[5:0] T606;
  wire[5:0] T607;
  wire[5:0] T608;
  wire[5:0] T609;
  wire[5:0] T610;
  wire[5:0] T611;
  wire[5:0] T612;
  wire[5:0] T613;
  wire[5:0] T614;
  wire[5:0] T615;
  wire T616;
  wire[54:0] T11;
  wire[22:0] T12;
  wire[6:0] T13;
  wire[2:0] T14;
  wire T15;
  wire[2:0] T16;
  wire[6:0] T17;
  wire[22:0] T18;
  wire[54:0] notCDom_reduced2AbsSigSum;
  wire[54:0] T19;
  wire[27:0] T20;
  wire[13:0] T21;
  wire[6:0] T22;
  wire[3:0] T23;
  wire[1:0] T24;
  wire T25;
  wire T26;
  wire[1:0] T27;
  wire[108:0] notCDom_absSigSum;
  wire[108:0] T28;
  wire[108:0] T617;
  wire[108:0] T29;
  wire[161:0] sigSum;
  wire[106:0] T30;
  wire[105:0] T31;
  wire[54:0] T32;
  wire[54:0] T33;
  wire T34;
  wire[108:0] T35;
  wire[108:0] T36;
  wire notCDom_signSigSum;
  wire T37;
  wire T38;
  wire[1:0] T39;
  wire[1:0] T40;
  wire T41;
  wire T42;
  wire[1:0] T43;
  wire T44;
  wire T45;
  wire[1:0] T46;
  wire[2:0] T47;
  wire[1:0] T48;
  wire T49;
  wire T50;
  wire[1:0] T51;
  wire T52;
  wire T53;
  wire[1:0] T54;
  wire T55;
  wire T56;
  wire[1:0] T57;
  wire[6:0] T58;
  wire[3:0] T59;
  wire[1:0] T60;
  wire T61;
  wire T62;
  wire[1:0] T63;
  wire T64;
  wire T65;
  wire[1:0] T66;
  wire[1:0] T67;
  wire T68;
  wire T69;
  wire[1:0] T70;
  wire T71;
  wire T72;
  wire[1:0] T73;
  wire[2:0] T74;
  wire[1:0] T75;
  wire T76;
  wire T77;
  wire[1:0] T78;
  wire T79;
  wire T80;
  wire[1:0] T81;
  wire T82;
  wire T83;
  wire[1:0] T84;
  wire[13:0] T85;
  wire[6:0] T86;
  wire[3:0] T87;
  wire[1:0] T88;
  wire T89;
  wire T90;
  wire[1:0] T91;
  wire T92;
  wire T93;
  wire[1:0] T94;
  wire[1:0] T95;
  wire T96;
  wire T97;
  wire[1:0] T98;
  wire T99;
  wire T100;
  wire[1:0] T101;
  wire[2:0] T102;
  wire[1:0] T103;
  wire T104;
  wire T105;
  wire[1:0] T106;
  wire T107;
  wire T108;
  wire[1:0] T109;
  wire T110;
  wire T111;
  wire[1:0] T112;
  wire[6:0] T113;
  wire[3:0] T114;
  wire[1:0] T115;
  wire T116;
  wire T117;
  wire[1:0] T118;
  wire T119;
  wire T120;
  wire[1:0] T121;
  wire[1:0] T122;
  wire T123;
  wire T124;
  wire[1:0] T125;
  wire T126;
  wire T127;
  wire[1:0] T128;
  wire[2:0] T129;
  wire[1:0] T130;
  wire T131;
  wire T132;
  wire[1:0] T133;
  wire T134;
  wire T135;
  wire[1:0] T136;
  wire T137;
  wire T138;
  wire[1:0] T139;
  wire[26:0] T140;
  wire[13:0] T141;
  wire[6:0] T142;
  wire[3:0] T143;
  wire[1:0] T144;
  wire T145;
  wire T146;
  wire[1:0] T147;
  wire T148;
  wire T149;
  wire[1:0] T150;
  wire[1:0] T151;
  wire T152;
  wire T153;
  wire[1:0] T154;
  wire T155;
  wire T156;
  wire[1:0] T157;
  wire[2:0] T158;
  wire[1:0] T159;
  wire T160;
  wire T161;
  wire[1:0] T162;
  wire T163;
  wire T164;
  wire[1:0] T165;
  wire T166;
  wire T167;
  wire[1:0] T168;
  wire[6:0] T169;
  wire[3:0] T170;
  wire[1:0] T171;
  wire T172;
  wire T173;
  wire[1:0] T174;
  wire T175;
  wire T176;
  wire[1:0] T177;
  wire[1:0] T178;
  wire T179;
  wire T180;
  wire[1:0] T181;
  wire T182;
  wire T183;
  wire[1:0] T184;
  wire[2:0] T185;
  wire[1:0] T186;
  wire T187;
  wire T188;
  wire[1:0] T189;
  wire T190;
  wire T191;
  wire[1:0] T192;
  wire T193;
  wire T194;
  wire[1:0] T195;
  wire[12:0] T196;
  wire[6:0] T197;
  wire[3:0] T198;
  wire[1:0] T199;
  wire T200;
  wire T201;
  wire[1:0] T202;
  wire T203;
  wire T204;
  wire[1:0] T205;
  wire[1:0] T206;
  wire T207;
  wire T208;
  wire[1:0] T209;
  wire T210;
  wire T211;
  wire[1:0] T212;
  wire[2:0] T213;
  wire[1:0] T214;
  wire T215;
  wire T216;
  wire[1:0] T217;
  wire T218;
  wire T219;
  wire[1:0] T220;
  wire T221;
  wire T222;
  wire[1:0] T223;
  wire[5:0] T224;
  wire[2:0] T225;
  wire[1:0] T226;
  wire T227;
  wire T228;
  wire[1:0] T229;
  wire T230;
  wire T231;
  wire[1:0] T232;
  wire T233;
  wire T234;
  wire[1:0] T235;
  wire[2:0] T236;
  wire[1:0] T237;
  wire T238;
  wire T239;
  wire[1:0] T240;
  wire T241;
  wire T242;
  wire[1:0] T243;
  wire T244;
  wire T245;
  wire T246;
  wire[1:0] T247;
  wire T248;
  wire[1:0] T249;
  wire T250;
  wire[3:0] T251;
  wire[1:0] T252;
  wire T253;
  wire[1:0] T254;
  wire[3:0] T255;
  wire T256;
  wire[1:0] T257;
  wire T258;
  wire[1:0] T259;
  wire T260;
  wire[15:0] T261;
  wire[15:0] T262;
  wire[15:0] T263;
  wire[14:0] T264;
  wire[15:0] T265;
  wire[15:0] T266;
  wire[15:0] T267;
  wire[13:0] T268;
  wire[15:0] T269;
  wire[15:0] T270;
  wire[15:0] T271;
  wire[11:0] T272;
  wire[15:0] T273;
  wire[15:0] T274;
  wire[15:0] T275;
  wire[7:0] T276;
  wire[15:0] T277;
  wire[15:0] T278;
  wire[15:0] T618;
  wire[7:0] T279;
  wire[15:0] T280;
  wire[15:0] T619;
  wire[11:0] T281;
  wire[15:0] T282;
  wire[15:0] T620;
  wire[13:0] T283;
  wire[15:0] T284;
  wire[15:0] T621;
  wire[14:0] T285;
  wire[31:0] T286;
  wire[31:0] T287;
  wire[31:0] T288;
  wire[30:0] T289;
  wire[31:0] T290;
  wire[31:0] T291;
  wire[31:0] T292;
  wire[29:0] T293;
  wire[31:0] T294;
  wire[31:0] T295;
  wire[31:0] T296;
  wire[27:0] T297;
  wire[31:0] T298;
  wire[31:0] T299;
  wire[31:0] T300;
  wire[23:0] T301;
  wire[31:0] T302;
  wire[31:0] T303;
  wire[31:0] T304;
  wire[15:0] T305;
  wire[31:0] T306;
  wire[31:0] T307;
  wire[31:0] T622;
  wire[15:0] T308;
  wire[31:0] T309;
  wire[31:0] T623;
  wire[23:0] T310;
  wire[31:0] T311;
  wire[31:0] T624;
  wire[27:0] T312;
  wire[31:0] T313;
  wire[31:0] T625;
  wire[29:0] T314;
  wire[31:0] T315;
  wire[31:0] T626;
  wire[30:0] T316;
  wire T627;
  wire T628;
  wire T629;
  wire T630;
  wire T631;
  wire T632;
  wire T633;
  wire T634;
  wire T635;
  wire T636;
  wire T637;
  wire T638;
  wire T639;
  wire T640;
  wire T641;
  wire T642;
  wire T643;
  wire T644;
  wire T645;
  wire T646;
  wire T647;
  wire T648;
  wire T649;
  wire T650;
  wire T651;
  wire T652;
  wire T653;
  wire T654;
  wire T655;
  wire T656;
  wire T657;
  wire T658;
  wire T659;
  wire T660;
  wire T661;
  wire T662;
  wire T663;
  wire T664;
  wire T665;
  wire T666;
  wire T667;
  wire T668;
  wire T669;
  wire T670;
  wire T671;
  wire T672;
  wire T673;
  wire T674;
  wire T675;
  wire T676;
  wire T677;
  wire T678;
  wire T679;
  wire[3:0] T317;
  wire[1:0] T318;
  wire T319;
  wire[1:0] T320;
  wire[3:0] T321;
  wire T322;
  wire[1:0] T323;
  wire T324;
  wire[1:0] T325;
  wire T326;
  wire[7:0] T327;
  wire[7:0] T328;
  wire[7:0] T329;
  wire[6:0] T330;
  wire[7:0] T331;
  wire[7:0] T332;
  wire[7:0] T333;
  wire[5:0] T334;
  wire[7:0] T335;
  wire[7:0] T336;
  wire[7:0] T337;
  wire[3:0] T338;
  wire[7:0] T339;
  wire[7:0] T340;
  wire[7:0] T680;
  wire[3:0] T341;
  wire[7:0] T342;
  wire[7:0] T681;
  wire[5:0] T343;
  wire[7:0] T344;
  wire[7:0] T682;
  wire[6:0] T345;
  wire[13:0] T346;
  wire[13:0] T347;
  wire[6:0] T348;
  wire[3:0] T349;
  wire[1:0] T350;
  wire T351;
  wire T352;
  wire[1:0] T353;
  wire[26:0] T354;
  wire[26:0] T355;
  wire T356;
  wire T357;
  wire[1:0] T358;
  wire[1:0] T359;
  wire T360;
  wire T361;
  wire[1:0] T362;
  wire T363;
  wire T364;
  wire[1:0] T365;
  wire[2:0] T366;
  wire[1:0] T367;
  wire T368;
  wire T369;
  wire[1:0] T370;
  wire T371;
  wire T372;
  wire[1:0] T373;
  wire T374;
  wire T375;
  wire[1:0] T376;
  wire[6:0] T377;
  wire[3:0] T378;
  wire[1:0] T379;
  wire T380;
  wire T381;
  wire[1:0] T382;
  wire T383;
  wire T384;
  wire[1:0] T385;
  wire[1:0] T386;
  wire T387;
  wire T388;
  wire[1:0] T389;
  wire T390;
  wire T391;
  wire[1:0] T392;
  wire[2:0] T393;
  wire[1:0] T394;
  wire T395;
  wire T396;
  wire[1:0] T397;
  wire T398;
  wire T399;
  wire[1:0] T400;
  wire T401;
  wire T402;
  wire T403;
  wire T404;
  wire[2:0] T405;
  wire[57:0] notCDom_mainSig;
  wire[235:0] T406;
  wire[6:0] notCDom_nearNormDist;
  wire[54:0] T407;
  wire[55:0] CDom_sig;
  wire T408;
  wire CDom_absSigSumExtra;
  wire T409;
  wire[53:0] T410;
  wire T411;
  wire[52:0] T412;
  wire[52:0] T413;
  wire T414;
  wire CDom_reduced4SigExtra;
  wire[13:0] T415;
  wire[13:0] T683;
  wire[12:0] T416;
  wire[4:0] T417;
  wire T418;
  wire[4:0] T419;
  wire[12:0] T420;
  wire[16:0] T421;
  wire[3:0] T422;
  wire[3:0] T423;
  wire[3:0] T424;
  wire[1:0] T425;
  wire T426;
  wire[1:0] T427;
  wire[3:0] T428;
  wire T429;
  wire[1:0] T430;
  wire T431;
  wire[1:0] T432;
  wire T433;
  wire[7:0] T434;
  wire[7:0] T435;
  wire[7:0] T436;
  wire[6:0] T437;
  wire[7:0] T438;
  wire[7:0] T439;
  wire[7:0] T440;
  wire[5:0] T441;
  wire[7:0] T442;
  wire[7:0] T443;
  wire[7:0] T444;
  wire[3:0] T445;
  wire[7:0] T446;
  wire[7:0] T447;
  wire[7:0] T684;
  wire[3:0] T448;
  wire[7:0] T449;
  wire[7:0] T685;
  wire[5:0] T450;
  wire[7:0] T451;
  wire[7:0] T686;
  wire[6:0] T452;
  wire[13:0] T453;
  wire[13:0] T454;
  wire[6:0] T455;
  wire[3:0] T456;
  wire[1:0] T457;
  wire T458;
  wire T459;
  wire[3:0] T460;
  wire[54:0] T461;
  wire[52:0] T462;
  wire[107:0] CDom_absSigSum;
  wire[107:0] T463;
  wire[106:0] T464;
  wire[104:0] T465;
  wire[1:0] T466;
  wire[107:0] T467;
  wire[107:0] T468;
  wire T469;
  wire T470;
  wire[3:0] T471;
  wire[1:0] T472;
  wire T473;
  wire T474;
  wire[3:0] T475;
  wire T476;
  wire T477;
  wire[3:0] T478;
  wire[2:0] T479;
  wire[1:0] T480;
  wire T481;
  wire T482;
  wire[3:0] T483;
  wire T484;
  wire T485;
  wire[3:0] T486;
  wire T487;
  wire T488;
  wire[3:0] T489;
  wire[6:0] T490;
  wire[3:0] T491;
  wire[1:0] T492;
  wire T493;
  wire T494;
  wire[3:0] T495;
  wire T496;
  wire T497;
  wire[3:0] T498;
  wire[1:0] T499;
  wire T500;
  wire T501;
  wire[3:0] T502;
  wire T503;
  wire T504;
  wire[3:0] T505;
  wire[2:0] T506;
  wire[1:0] T507;
  wire T508;
  wire T509;
  wire[3:0] T510;
  wire T511;
  wire T512;
  wire[3:0] T513;
  wire T514;
  wire T515;
  wire[2:0] T516;
  wire T517;
  wire[2:0] T518;
  wire[57:0] CDom_mainSig;
  wire[170:0] T519;
  wire[54:0] T520;
  wire[12:0] T521;
  wire[12:0] notCDom_sExp;
  wire[12:0] T687;
  wire[7:0] T522;
  wire[7:0] T523;
  wire[4:0] T688;
  wire T689;
  wire[12:0] CDom_sExp;
  wire[12:0] T690;
  wire[1:0] T524;
  wire[1:0] T525;
  wire[10:0] T691;
  wire T692;
  wire T526;
  wire T527;
  wire T528;
  wire notCDom_sign;
  wire T529;
  wire roundingMode_min;
  wire notCDom_completeCancellation;
  wire[1:0] T530;
  wire CDom_sign;
  wire T531;
  wire T532;
  wire notNaN_addZeros;
  wire T533;
  wire T534;
  wire notNaN_isInfOut;
  wire notNaN_isInfProd;
  wire T535;
  wire T536;
  wire T537;
  wire T538;
  wire T539;
  wire T540;
  wire T541;
  wire T542;
  wire T543;
  wire T544;
  wire T545;
  wire T546;
  wire T547;
  wire T548;
  wire T549;
  wire T550;
  wire T551;
  wire T552;
  wire T553;
  wire T554;
  wire T555;
  wire T556;
  wire T557;
  wire T558;
  wire T559;
  wire T560;


  assign io_rawOut_sig = T0;
  assign T0 = io_fromPreMul_CIsDominant ? CDom_sig : notCDom_sig;
  assign notCDom_sig = {T407, T1};
  assign T1 = T404 | notCDom_reduced4SigExtra;
  assign notCDom_reduced4SigExtra = T2 != 14'h0;
  assign T2 = T346 & T561;
  assign T561 = {1'h0, T3};
  assign T3 = {T327, T4};
  assign T4 = {T317, T5};
  assign T5 = T6[4];
  assign T6 = T7[12:8];
  assign T7 = T8[13:1];
  assign T8 = $signed(33'h100000000) >>> T9;
  assign T9 = ~ T10;
  assign T10 = T562 >> 1'h1;
  assign T562 = T679 ? 1'h0 : T563;
  assign T563 = T678 ? 1'h1 : T564;
  assign T564 = T677 ? 2'h2 : T565;
  assign T565 = T676 ? 2'h3 : T566;
  assign T566 = T675 ? 3'h4 : T567;
  assign T567 = T674 ? 3'h5 : T568;
  assign T568 = T673 ? 3'h6 : T569;
  assign T569 = T672 ? 3'h7 : T570;
  assign T570 = T671 ? 4'h8 : T571;
  assign T571 = T670 ? 4'h9 : T572;
  assign T572 = T669 ? 4'ha : T573;
  assign T573 = T668 ? 4'hb : T574;
  assign T574 = T667 ? 4'hc : T575;
  assign T575 = T666 ? 4'hd : T576;
  assign T576 = T665 ? 4'he : T577;
  assign T577 = T664 ? 4'hf : T578;
  assign T578 = T663 ? 5'h10 : T579;
  assign T579 = T662 ? 5'h11 : T580;
  assign T580 = T661 ? 5'h12 : T581;
  assign T581 = T660 ? 5'h13 : T582;
  assign T582 = T659 ? 5'h14 : T583;
  assign T583 = T658 ? 5'h15 : T584;
  assign T584 = T657 ? 5'h16 : T585;
  assign T585 = T656 ? 5'h17 : T586;
  assign T586 = T655 ? 5'h18 : T587;
  assign T587 = T654 ? 5'h19 : T588;
  assign T588 = T653 ? 5'h1a : T589;
  assign T589 = T652 ? 5'h1b : T590;
  assign T590 = T651 ? 5'h1c : T591;
  assign T591 = T650 ? 5'h1d : T592;
  assign T592 = T649 ? 5'h1e : T593;
  assign T593 = T648 ? 5'h1f : T594;
  assign T594 = T647 ? 6'h20 : T595;
  assign T595 = T646 ? 6'h21 : T596;
  assign T596 = T645 ? 6'h22 : T597;
  assign T597 = T644 ? 6'h23 : T598;
  assign T598 = T643 ? 6'h24 : T599;
  assign T599 = T642 ? 6'h25 : T600;
  assign T600 = T641 ? 6'h26 : T601;
  assign T601 = T640 ? 6'h27 : T602;
  assign T602 = T639 ? 6'h28 : T603;
  assign T603 = T638 ? 6'h29 : T604;
  assign T604 = T637 ? 6'h2a : T605;
  assign T605 = T636 ? 6'h2b : T606;
  assign T606 = T635 ? 6'h2c : T607;
  assign T607 = T634 ? 6'h2d : T608;
  assign T608 = T633 ? 6'h2e : T609;
  assign T609 = T632 ? 6'h2f : T610;
  assign T610 = T631 ? 6'h30 : T611;
  assign T611 = T630 ? 6'h31 : T612;
  assign T612 = T629 ? 6'h32 : T613;
  assign T613 = T628 ? 6'h33 : T614;
  assign T614 = T627 ? 6'h34 : T615;
  assign T615 = T616 ? 6'h35 : 6'h36;
  assign T616 = T11[53];
  assign T11 = {T286, T12};
  assign T12 = {T261, T13};
  assign T13 = {T251, T14};
  assign T14 = {T247, T15};
  assign T15 = T16[2];
  assign T16 = T17[6:4];
  assign T17 = T18[22:16];
  assign T18 = notCDom_reduced2AbsSigSum[54:32];
  assign notCDom_reduced2AbsSigSum = T19;
  assign T19 = {T140, T20};
  assign T20 = {T85, T21};
  assign T21 = {T58, T22};
  assign T22 = {T47, T23};
  assign T23 = {T40, T24};
  assign T24 = {T37, T25};
  assign T25 = T26;
  assign T26 = T27 != 2'h0;
  assign T27 = notCDom_absSigSum[1:0];
  assign notCDom_absSigSum = notCDom_signSigSum ? T35 : T28;
  assign T28 = T29 + T617;
  assign T617 = {108'h0, io_fromPreMul_doSubMags};
  assign T29 = sigSum[108:0];
  assign sigSum = {T32, T30};
  assign T30 = {T31, io_fromPreMul_bit0AlignedSigC};
  assign T31 = io_mulAddResult[105:0];
  assign T32 = T34 ? T33 : io_fromPreMul_highAlignedSigC;
  assign T33 = io_fromPreMul_highAlignedSigC + 55'h1;
  assign T34 = io_mulAddResult[106];
  assign T35 = ~ T36;
  assign T36 = sigSum[108:0];
  assign notCDom_signSigSum = sigSum[109];
  assign T37 = T38;
  assign T38 = T39 != 2'h0;
  assign T39 = notCDom_absSigSum[3:2];
  assign T40 = {T44, T41};
  assign T41 = T42;
  assign T42 = T43 != 2'h0;
  assign T43 = notCDom_absSigSum[5:4];
  assign T44 = T45;
  assign T45 = T46 != 2'h0;
  assign T46 = notCDom_absSigSum[7:6];
  assign T47 = {T55, T48};
  assign T48 = {T52, T49};
  assign T49 = T50;
  assign T50 = T51 != 2'h0;
  assign T51 = notCDom_absSigSum[9:8];
  assign T52 = T53;
  assign T53 = T54 != 2'h0;
  assign T54 = notCDom_absSigSum[11:10];
  assign T55 = T56;
  assign T56 = T57 != 2'h0;
  assign T57 = notCDom_absSigSum[13:12];
  assign T58 = {T74, T59};
  assign T59 = {T67, T60};
  assign T60 = {T64, T61};
  assign T61 = T62;
  assign T62 = T63 != 2'h0;
  assign T63 = notCDom_absSigSum[15:14];
  assign T64 = T65;
  assign T65 = T66 != 2'h0;
  assign T66 = notCDom_absSigSum[17:16];
  assign T67 = {T71, T68};
  assign T68 = T69;
  assign T69 = T70 != 2'h0;
  assign T70 = notCDom_absSigSum[19:18];
  assign T71 = T72;
  assign T72 = T73 != 2'h0;
  assign T73 = notCDom_absSigSum[21:20];
  assign T74 = {T82, T75};
  assign T75 = {T79, T76};
  assign T76 = T77;
  assign T77 = T78 != 2'h0;
  assign T78 = notCDom_absSigSum[23:22];
  assign T79 = T80;
  assign T80 = T81 != 2'h0;
  assign T81 = notCDom_absSigSum[25:24];
  assign T82 = T83;
  assign T83 = T84 != 2'h0;
  assign T84 = notCDom_absSigSum[27:26];
  assign T85 = {T113, T86};
  assign T86 = {T102, T87};
  assign T87 = {T95, T88};
  assign T88 = {T92, T89};
  assign T89 = T90;
  assign T90 = T91 != 2'h0;
  assign T91 = notCDom_absSigSum[29:28];
  assign T92 = T93;
  assign T93 = T94 != 2'h0;
  assign T94 = notCDom_absSigSum[31:30];
  assign T95 = {T99, T96};
  assign T96 = T97;
  assign T97 = T98 != 2'h0;
  assign T98 = notCDom_absSigSum[33:32];
  assign T99 = T100;
  assign T100 = T101 != 2'h0;
  assign T101 = notCDom_absSigSum[35:34];
  assign T102 = {T110, T103};
  assign T103 = {T107, T104};
  assign T104 = T105;
  assign T105 = T106 != 2'h0;
  assign T106 = notCDom_absSigSum[37:36];
  assign T107 = T108;
  assign T108 = T109 != 2'h0;
  assign T109 = notCDom_absSigSum[39:38];
  assign T110 = T111;
  assign T111 = T112 != 2'h0;
  assign T112 = notCDom_absSigSum[41:40];
  assign T113 = {T129, T114};
  assign T114 = {T122, T115};
  assign T115 = {T119, T116};
  assign T116 = T117;
  assign T117 = T118 != 2'h0;
  assign T118 = notCDom_absSigSum[43:42];
  assign T119 = T120;
  assign T120 = T121 != 2'h0;
  assign T121 = notCDom_absSigSum[45:44];
  assign T122 = {T126, T123};
  assign T123 = T124;
  assign T124 = T125 != 2'h0;
  assign T125 = notCDom_absSigSum[47:46];
  assign T126 = T127;
  assign T127 = T128 != 2'h0;
  assign T128 = notCDom_absSigSum[49:48];
  assign T129 = {T137, T130};
  assign T130 = {T134, T131};
  assign T131 = T132;
  assign T132 = T133 != 2'h0;
  assign T133 = notCDom_absSigSum[51:50];
  assign T134 = T135;
  assign T135 = T136 != 2'h0;
  assign T136 = notCDom_absSigSum[53:52];
  assign T137 = T138;
  assign T138 = T139 != 2'h0;
  assign T139 = notCDom_absSigSum[55:54];
  assign T140 = {T196, T141};
  assign T141 = {T169, T142};
  assign T142 = {T158, T143};
  assign T143 = {T151, T144};
  assign T144 = {T148, T145};
  assign T145 = T146;
  assign T146 = T147 != 2'h0;
  assign T147 = notCDom_absSigSum[57:56];
  assign T148 = T149;
  assign T149 = T150 != 2'h0;
  assign T150 = notCDom_absSigSum[59:58];
  assign T151 = {T155, T152};
  assign T152 = T153;
  assign T153 = T154 != 2'h0;
  assign T154 = notCDom_absSigSum[61:60];
  assign T155 = T156;
  assign T156 = T157 != 2'h0;
  assign T157 = notCDom_absSigSum[63:62];
  assign T158 = {T166, T159};
  assign T159 = {T163, T160};
  assign T160 = T161;
  assign T161 = T162 != 2'h0;
  assign T162 = notCDom_absSigSum[65:64];
  assign T163 = T164;
  assign T164 = T165 != 2'h0;
  assign T165 = notCDom_absSigSum[67:66];
  assign T166 = T167;
  assign T167 = T168 != 2'h0;
  assign T168 = notCDom_absSigSum[69:68];
  assign T169 = {T185, T170};
  assign T170 = {T178, T171};
  assign T171 = {T175, T172};
  assign T172 = T173;
  assign T173 = T174 != 2'h0;
  assign T174 = notCDom_absSigSum[71:70];
  assign T175 = T176;
  assign T176 = T177 != 2'h0;
  assign T177 = notCDom_absSigSum[73:72];
  assign T178 = {T182, T179};
  assign T179 = T180;
  assign T180 = T181 != 2'h0;
  assign T181 = notCDom_absSigSum[75:74];
  assign T182 = T183;
  assign T183 = T184 != 2'h0;
  assign T184 = notCDom_absSigSum[77:76];
  assign T185 = {T193, T186};
  assign T186 = {T190, T187};
  assign T187 = T188;
  assign T188 = T189 != 2'h0;
  assign T189 = notCDom_absSigSum[79:78];
  assign T190 = T191;
  assign T191 = T192 != 2'h0;
  assign T192 = notCDom_absSigSum[81:80];
  assign T193 = T194;
  assign T194 = T195 != 2'h0;
  assign T195 = notCDom_absSigSum[83:82];
  assign T196 = {T224, T197};
  assign T197 = {T213, T198};
  assign T198 = {T206, T199};
  assign T199 = {T203, T200};
  assign T200 = T201;
  assign T201 = T202 != 2'h0;
  assign T202 = notCDom_absSigSum[85:84];
  assign T203 = T204;
  assign T204 = T205 != 2'h0;
  assign T205 = notCDom_absSigSum[87:86];
  assign T206 = {T210, T207};
  assign T207 = T208;
  assign T208 = T209 != 2'h0;
  assign T209 = notCDom_absSigSum[89:88];
  assign T210 = T211;
  assign T211 = T212 != 2'h0;
  assign T212 = notCDom_absSigSum[91:90];
  assign T213 = {T221, T214};
  assign T214 = {T218, T215};
  assign T215 = T216;
  assign T216 = T217 != 2'h0;
  assign T217 = notCDom_absSigSum[93:92];
  assign T218 = T219;
  assign T219 = T220 != 2'h0;
  assign T220 = notCDom_absSigSum[95:94];
  assign T221 = T222;
  assign T222 = T223 != 2'h0;
  assign T223 = notCDom_absSigSum[97:96];
  assign T224 = {T236, T225};
  assign T225 = {T233, T226};
  assign T226 = {T230, T227};
  assign T227 = T228;
  assign T228 = T229 != 2'h0;
  assign T229 = notCDom_absSigSum[99:98];
  assign T230 = T231;
  assign T231 = T232 != 2'h0;
  assign T232 = notCDom_absSigSum[101:100];
  assign T233 = T234;
  assign T234 = T235 != 2'h0;
  assign T235 = notCDom_absSigSum[103:102];
  assign T236 = {T244, T237};
  assign T237 = {T241, T238};
  assign T238 = T239;
  assign T239 = T240 != 2'h0;
  assign T240 = notCDom_absSigSum[105:104];
  assign T241 = T242;
  assign T242 = T243 != 2'h0;
  assign T243 = notCDom_absSigSum[107:106];
  assign T244 = T245;
  assign T245 = T246 != 1'h0;
  assign T246 = notCDom_absSigSum[108];
  assign T247 = {T250, T248};
  assign T248 = T249[1];
  assign T249 = T16[1:0];
  assign T250 = T249[0];
  assign T251 = {T257, T252};
  assign T252 = {T256, T253};
  assign T253 = T254[1];
  assign T254 = T255[3:2];
  assign T255 = T17[3:0];
  assign T256 = T254[0];
  assign T257 = {T260, T258};
  assign T258 = T259[1];
  assign T259 = T255[1:0];
  assign T260 = T259[0];
  assign T261 = T284 | T262;
  assign T262 = T263 & 16'haaaa;
  assign T263 = T264 << 1'h1;
  assign T264 = T265[14:0];
  assign T265 = T282 | T266;
  assign T266 = T267 & 16'hcccc;
  assign T267 = T268 << 2'h2;
  assign T268 = T269[13:0];
  assign T269 = T280 | T270;
  assign T270 = T271 & 16'hf0f0;
  assign T271 = T272 << 3'h4;
  assign T272 = T273[11:0];
  assign T273 = T278 | T274;
  assign T274 = T275 & 16'hff00;
  assign T275 = T276 << 4'h8;
  assign T276 = T277[7:0];
  assign T277 = T18[15:0];
  assign T278 = T618 & 16'hff;
  assign T618 = {8'h0, T279};
  assign T279 = T277 >> 4'h8;
  assign T280 = T619 & 16'hf0f;
  assign T619 = {4'h0, T281};
  assign T281 = T273 >> 3'h4;
  assign T282 = T620 & 16'h3333;
  assign T620 = {2'h0, T283};
  assign T283 = T269 >> 2'h2;
  assign T284 = T621 & 16'h5555;
  assign T621 = {1'h0, T285};
  assign T285 = T265 >> 1'h1;
  assign T286 = T315 | T287;
  assign T287 = T288 & 32'haaaaaaaa;
  assign T288 = T289 << 1'h1;
  assign T289 = T290[30:0];
  assign T290 = T313 | T291;
  assign T291 = T292 & 32'hcccccccc;
  assign T292 = T293 << 2'h2;
  assign T293 = T294[29:0];
  assign T294 = T311 | T295;
  assign T295 = T296 & 32'hf0f0f0f0;
  assign T296 = T297 << 3'h4;
  assign T297 = T298[27:0];
  assign T298 = T309 | T299;
  assign T299 = T300 & 32'hff00ff00;
  assign T300 = T301 << 4'h8;
  assign T301 = T302[23:0];
  assign T302 = T307 | T303;
  assign T303 = T304 & 32'hffff0000;
  assign T304 = T305 << 5'h10;
  assign T305 = T306[15:0];
  assign T306 = notCDom_reduced2AbsSigSum[31:0];
  assign T307 = T622 & 32'hffff;
  assign T622 = {16'h0, T308};
  assign T308 = T306 >> 5'h10;
  assign T309 = T623 & 32'hff00ff;
  assign T623 = {8'h0, T310};
  assign T310 = T302 >> 4'h8;
  assign T311 = T624 & 32'hf0f0f0f;
  assign T624 = {4'h0, T312};
  assign T312 = T298 >> 3'h4;
  assign T313 = T625 & 32'h33333333;
  assign T625 = {2'h0, T314};
  assign T314 = T294 >> 2'h2;
  assign T315 = T626 & 32'h55555555;
  assign T626 = {1'h0, T316};
  assign T316 = T290 >> 1'h1;
  assign T627 = T11[52];
  assign T628 = T11[51];
  assign T629 = T11[50];
  assign T630 = T11[49];
  assign T631 = T11[48];
  assign T632 = T11[47];
  assign T633 = T11[46];
  assign T634 = T11[45];
  assign T635 = T11[44];
  assign T636 = T11[43];
  assign T637 = T11[42];
  assign T638 = T11[41];
  assign T639 = T11[40];
  assign T640 = T11[39];
  assign T641 = T11[38];
  assign T642 = T11[37];
  assign T643 = T11[36];
  assign T644 = T11[35];
  assign T645 = T11[34];
  assign T646 = T11[33];
  assign T647 = T11[32];
  assign T648 = T11[31];
  assign T649 = T11[30];
  assign T650 = T11[29];
  assign T651 = T11[28];
  assign T652 = T11[27];
  assign T653 = T11[26];
  assign T654 = T11[25];
  assign T655 = T11[24];
  assign T656 = T11[23];
  assign T657 = T11[22];
  assign T658 = T11[21];
  assign T659 = T11[20];
  assign T660 = T11[19];
  assign T661 = T11[18];
  assign T662 = T11[17];
  assign T663 = T11[16];
  assign T664 = T11[15];
  assign T665 = T11[14];
  assign T666 = T11[13];
  assign T667 = T11[12];
  assign T668 = T11[11];
  assign T669 = T11[10];
  assign T670 = T11[9];
  assign T671 = T11[8];
  assign T672 = T11[7];
  assign T673 = T11[6];
  assign T674 = T11[5];
  assign T675 = T11[4];
  assign T676 = T11[3];
  assign T677 = T11[2];
  assign T678 = T11[1];
  assign T679 = T11[0];
  assign T317 = {T323, T318};
  assign T318 = {T322, T319};
  assign T319 = T320[1];
  assign T320 = T321[3:2];
  assign T321 = T6[3:0];
  assign T322 = T320[0];
  assign T323 = {T326, T324};
  assign T324 = T325[1];
  assign T325 = T321[1:0];
  assign T326 = T325[0];
  assign T327 = T344 | T328;
  assign T328 = T329 & 8'haa;
  assign T329 = T330 << 1'h1;
  assign T330 = T331[6:0];
  assign T331 = T342 | T332;
  assign T332 = T333 & 8'hcc;
  assign T333 = T334 << 2'h2;
  assign T334 = T335[5:0];
  assign T335 = T340 | T336;
  assign T336 = T337 & 8'hf0;
  assign T337 = T338 << 3'h4;
  assign T338 = T339[3:0];
  assign T339 = T7[7:0];
  assign T340 = T680 & 8'hf;
  assign T680 = {4'h0, T341};
  assign T341 = T339 >> 3'h4;
  assign T342 = T681 & 8'h33;
  assign T681 = {2'h0, T343};
  assign T343 = T335 >> 2'h2;
  assign T344 = T682 & 8'h55;
  assign T682 = {1'h0, T345};
  assign T345 = T331 >> 1'h1;
  assign T346 = T347;
  assign T347 = {T377, T348};
  assign T348 = {T366, T349};
  assign T349 = {T359, T350};
  assign T350 = {T356, T351};
  assign T351 = T352;
  assign T352 = T353 != 2'h0;
  assign T353 = T354[1:0];
  assign T354 = T355 << 1'h0;
  assign T355 = notCDom_reduced2AbsSigSum[26:0];
  assign T356 = T357;
  assign T357 = T358 != 2'h0;
  assign T358 = T354[3:2];
  assign T359 = {T363, T360};
  assign T360 = T361;
  assign T361 = T362 != 2'h0;
  assign T362 = T354[5:4];
  assign T363 = T364;
  assign T364 = T365 != 2'h0;
  assign T365 = T354[7:6];
  assign T366 = {T374, T367};
  assign T367 = {T371, T368};
  assign T368 = T369;
  assign T369 = T370 != 2'h0;
  assign T370 = T354[9:8];
  assign T371 = T372;
  assign T372 = T373 != 2'h0;
  assign T373 = T354[11:10];
  assign T374 = T375;
  assign T375 = T376 != 2'h0;
  assign T376 = T354[13:12];
  assign T377 = {T393, T378};
  assign T378 = {T386, T379};
  assign T379 = {T383, T380};
  assign T380 = T381;
  assign T381 = T382 != 2'h0;
  assign T382 = T354[15:14];
  assign T383 = T384;
  assign T384 = T385 != 2'h0;
  assign T385 = T354[17:16];
  assign T386 = {T390, T387};
  assign T387 = T388;
  assign T388 = T389 != 2'h0;
  assign T389 = T354[19:18];
  assign T390 = T391;
  assign T391 = T392 != 2'h0;
  assign T392 = T354[21:20];
  assign T393 = {T401, T394};
  assign T394 = {T398, T395};
  assign T395 = T396;
  assign T396 = T397 != 2'h0;
  assign T397 = T354[23:22];
  assign T398 = T399;
  assign T399 = T400 != 2'h0;
  assign T400 = T354[25:24];
  assign T401 = T402;
  assign T402 = T403 != 1'h0;
  assign T403 = T354[26];
  assign T404 = T405 != 3'h0;
  assign T405 = notCDom_mainSig[2:0];
  assign notCDom_mainSig = T406[109:52];
  assign T406 = notCDom_absSigSum << notCDom_nearNormDist;
  assign notCDom_nearNormDist = T562 << 1'h1;
  assign T407 = notCDom_mainSig >> 2'h3;
  assign CDom_sig = {T520, T408};
  assign T408 = T414 | CDom_absSigSumExtra;
  assign CDom_absSigSumExtra = io_fromPreMul_doSubMags ? T411 : T409;
  assign T409 = T410 != 54'h0;
  assign T410 = sigSum[54:1];
  assign T411 = T412 != 53'h0;
  assign T412 = ~ T413;
  assign T413 = sigSum[53:1];
  assign T414 = T517 | CDom_reduced4SigExtra;
  assign CDom_reduced4SigExtra = T415 != 14'h0;
  assign T415 = T453 & T683;
  assign T683 = {1'h0, T416};
  assign T416 = {T434, T417};
  assign T417 = {T424, T418};
  assign T418 = T419[4];
  assign T419 = T420[12:8];
  assign T420 = T421[13:1];
  assign T421 = $signed(17'h10000) >>> T422;
  assign T422 = ~ T423;
  assign T423 = io_fromPreMul_CDom_CAlignDist >> 2'h2;
  assign T424 = {T430, T425};
  assign T425 = {T429, T426};
  assign T426 = T427[1];
  assign T427 = T428[3:2];
  assign T428 = T419[3:0];
  assign T429 = T427[0];
  assign T430 = {T433, T431};
  assign T431 = T432[1];
  assign T432 = T428[1:0];
  assign T433 = T432[0];
  assign T434 = T451 | T435;
  assign T435 = T436 & 8'haa;
  assign T436 = T437 << 1'h1;
  assign T437 = T438[6:0];
  assign T438 = T449 | T439;
  assign T439 = T440 & 8'hcc;
  assign T440 = T441 << 2'h2;
  assign T441 = T442[5:0];
  assign T442 = T447 | T443;
  assign T443 = T444 & 8'hf0;
  assign T444 = T445 << 3'h4;
  assign T445 = T446[3:0];
  assign T446 = T420[7:0];
  assign T447 = T684 & 8'hf;
  assign T684 = {4'h0, T448};
  assign T448 = T446 >> 3'h4;
  assign T449 = T685 & 8'h33;
  assign T685 = {2'h0, T450};
  assign T450 = T442 >> 2'h2;
  assign T451 = T686 & 8'h55;
  assign T686 = {1'h0, T452};
  assign T452 = T438 >> 1'h1;
  assign T453 = T454;
  assign T454 = {T490, T455};
  assign T455 = {T479, T456};
  assign T456 = {T472, T457};
  assign T457 = {T469, T458};
  assign T458 = T459;
  assign T459 = T460 != 4'h0;
  assign T460 = T461[3:0];
  assign T461 = T462 << 2'h2;
  assign T462 = CDom_absSigSum[52:0];
  assign CDom_absSigSum = io_fromPreMul_doSubMags ? T467 : T463;
  assign T463 = {1'h0, T464};
  assign T464 = {T466, T465};
  assign T465 = sigSum[159:55];
  assign T466 = io_fromPreMul_highAlignedSigC[54:53];
  assign T467 = ~ T468;
  assign T468 = sigSum[161:54];
  assign T469 = T470;
  assign T470 = T471 != 4'h0;
  assign T471 = T461[7:4];
  assign T472 = {T476, T473};
  assign T473 = T474;
  assign T474 = T475 != 4'h0;
  assign T475 = T461[11:8];
  assign T476 = T477;
  assign T477 = T478 != 4'h0;
  assign T478 = T461[15:12];
  assign T479 = {T487, T480};
  assign T480 = {T484, T481};
  assign T481 = T482;
  assign T482 = T483 != 4'h0;
  assign T483 = T461[19:16];
  assign T484 = T485;
  assign T485 = T486 != 4'h0;
  assign T486 = T461[23:20];
  assign T487 = T488;
  assign T488 = T489 != 4'h0;
  assign T489 = T461[27:24];
  assign T490 = {T506, T491};
  assign T491 = {T499, T492};
  assign T492 = {T496, T493};
  assign T493 = T494;
  assign T494 = T495 != 4'h0;
  assign T495 = T461[31:28];
  assign T496 = T497;
  assign T497 = T498 != 4'h0;
  assign T498 = T461[35:32];
  assign T499 = {T503, T500};
  assign T500 = T501;
  assign T501 = T502 != 4'h0;
  assign T502 = T461[39:36];
  assign T503 = T504;
  assign T504 = T505 != 4'h0;
  assign T505 = T461[43:40];
  assign T506 = {T514, T507};
  assign T507 = {T511, T508};
  assign T508 = T509;
  assign T509 = T510 != 4'h0;
  assign T510 = T461[47:44];
  assign T511 = T512;
  assign T512 = T513 != 4'h0;
  assign T513 = T461[51:48];
  assign T514 = T515;
  assign T515 = T516 != 3'h0;
  assign T516 = T461[54:52];
  assign T517 = T518 != 3'h0;
  assign T518 = CDom_mainSig[2:0];
  assign CDom_mainSig = T519[107:50];
  assign T519 = CDom_absSigSum << io_fromPreMul_CDom_CAlignDist;
  assign T520 = CDom_mainSig >> 2'h3;
  assign io_rawOut_sExp = T521;
  assign T521 = io_fromPreMul_CIsDominant ? CDom_sExp : notCDom_sExp;
  assign notCDom_sExp = io_fromPreMul_sExpSum - T687;
  assign T687 = {T688, T522};
  assign T522 = T523;
  assign T523 = {1'h0, notCDom_nearNormDist};
  assign T688 = T689 ? 5'h1f : 5'h0;
  assign T689 = T522[7];
  assign CDom_sExp = io_fromPreMul_sExpSum - T690;
  assign T690 = {T691, T524};
  assign T524 = T525;
  assign T525 = {1'h0, io_fromPreMul_doSubMags};
  assign T691 = T692 ? 11'h7ff : 11'h0;
  assign T692 = T524[1];
  assign io_rawOut_sign = T526;
  assign T526 = T535 | T527;
  assign T527 = T531 & T528;
  assign T528 = io_fromPreMul_CIsDominant ? CDom_sign : notCDom_sign;
  assign notCDom_sign = notCDom_completeCancellation ? roundingMode_min : T529;
  assign T529 = io_fromPreMul_signProd ^ notCDom_signSigSum;
  assign roundingMode_min = io_roundingMode == 3'h2;
  assign notCDom_completeCancellation = T530 == 2'h0;
  assign T530 = notCDom_sig[55:54];
  assign CDom_sign = io_fromPreMul_signProd ^ io_fromPreMul_doSubMags;
  assign T531 = T534 & T532;
  assign T532 = notNaN_addZeros ^ 1'h1;
  assign notNaN_addZeros = T533 & io_fromPreMul_isZeroC;
  assign T533 = io_fromPreMul_isZeroA | io_fromPreMul_isZeroB;
  assign T534 = notNaN_isInfOut ^ 1'h1;
  assign notNaN_isInfOut = notNaN_isInfProd | io_fromPreMul_isInfC;
  assign notNaN_isInfProd = io_fromPreMul_isInfA | io_fromPreMul_isInfB;
  assign T535 = T539 | T536;
  assign T536 = T538 & T537;
  assign T537 = io_fromPreMul_signProd | CDom_sign;
  assign T538 = notNaN_addZeros & roundingMode_min;
  assign T539 = T544 | T540;
  assign T540 = T541 & CDom_sign;
  assign T541 = T542 & io_fromPreMul_signProd;
  assign T542 = notNaN_addZeros & T543;
  assign T543 = roundingMode_min ^ 1'h1;
  assign T544 = T546 | T545;
  assign T545 = io_fromPreMul_isInfC & CDom_sign;
  assign T546 = notNaN_isInfProd & io_fromPreMul_signProd;
  assign io_rawOut_isZero = T547;
  assign T547 = notNaN_addZeros | T548;
  assign T548 = T549 & notCDom_completeCancellation;
  assign T549 = io_fromPreMul_CIsDominant ^ 1'h1;
  assign io_rawOut_isInf = notNaN_isInfOut;
  assign io_rawOut_isNaN = T550;
  assign T550 = io_fromPreMul_isNaNAOrB | io_fromPreMul_isNaNC;
  assign io_invalidExc = T551;
  assign T551 = T557 | T552;
  assign T552 = T553 & io_fromPreMul_doSubMags;
  assign T553 = T554 & io_fromPreMul_isInfC;
  assign T554 = T556 & T555;
  assign T555 = io_fromPreMul_isInfA | io_fromPreMul_isInfB;
  assign T556 = io_fromPreMul_isNaNAOrB ^ 1'h1;
  assign T557 = T559 | T558;
  assign T558 = io_fromPreMul_isZeroA & io_fromPreMul_isInfB;
  assign T559 = io_fromPreMul_isSigNaNAny | T560;
  assign T560 = io_fromPreMul_isInfA & io_fromPreMul_isZeroB;
endmodule

module RoundAnyRawFNToRecFN(
    input  io_invalidExc,
    input  io_infiniteExc,
    input  io_in_isNaN,
    input  io_in_isInf,
    input  io_in_isZero,
    input  io_in_sign,
    input [12:0] io_in_sExp,
    input [55:0] io_in_sig,
    input [2:0] io_roundingMode,
    input  io_detectTininess,
    output[64:0] io_out,
    output[4:0] io_exceptionFlags
);

  wire[4:0] T0;
  wire[2:0] T1;
  wire[1:0] T2;
  wire inexact;
  wire T3;
  wire common_inexact;
  wire T4;
  wire T5;
  wire T6;
  wire[55:0] T7;
  wire[55:0] T8;
  wire[54:0] T9;
  wire[55:0] T10;
  wire[53:0] T11;
  wire[53:0] T240;
  wire doShiftSigDown1;
  wire[53:0] T12;
  wire[53:0] T13;
  wire[53:0] T241;
  wire[2:0] T14;
  wire[2:0] T15;
  wire[2:0] T16;
  wire[2:0] T17;
  wire[2:0] T18;
  wire T19;
  wire[2:0] T20;
  wire[64:0] T21;
  wire[5:0] T22;
  wire[6:0] T23;
  wire[7:0] T24;
  wire[8:0] T25;
  wire[9:0] T26;
  wire[10:0] T27;
  wire[11:0] T28;
  wire[11:0] T29;
  wire[1:0] T30;
  wire T31;
  wire[1:0] T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire[53:0] T38;
  wire[50:0] T39;
  wire[50:0] T40;
  wire[50:0] T41;
  wire[50:0] T42;
  wire[50:0] T43;
  wire[50:0] T44;
  wire[50:0] T45;
  wire[50:0] T46;
  wire[50:0] T47;
  wire[50:0] T48;
  wire[50:0] T49;
  wire[50:0] T50;
  wire[50:0] T51;
  wire[18:0] T52;
  wire[2:0] T53;
  wire T54;
  wire[2:0] T55;
  wire[18:0] T56;
  wire[50:0] T57;
  wire[64:0] T58;
  wire[5:0] T59;
  wire[6:0] T60;
  wire[7:0] T61;
  wire[8:0] T62;
  wire[1:0] T63;
  wire T64;
  wire[1:0] T65;
  wire T66;
  wire[15:0] T67;
  wire[15:0] T68;
  wire[15:0] T69;
  wire[14:0] T70;
  wire[15:0] T71;
  wire[15:0] T72;
  wire[15:0] T73;
  wire[13:0] T74;
  wire[15:0] T75;
  wire[15:0] T76;
  wire[15:0] T77;
  wire[11:0] T78;
  wire[15:0] T79;
  wire[15:0] T80;
  wire[15:0] T81;
  wire[7:0] T82;
  wire[15:0] T83;
  wire[15:0] T84;
  wire[15:0] T242;
  wire[7:0] T85;
  wire[15:0] T86;
  wire[15:0] T243;
  wire[11:0] T87;
  wire[15:0] T88;
  wire[15:0] T244;
  wire[13:0] T89;
  wire[15:0] T90;
  wire[15:0] T245;
  wire[14:0] T91;
  wire[31:0] T92;
  wire[31:0] T93;
  wire[31:0] T94;
  wire[30:0] T95;
  wire[31:0] T96;
  wire[31:0] T97;
  wire[31:0] T98;
  wire[29:0] T99;
  wire[31:0] T100;
  wire[31:0] T101;
  wire[31:0] T102;
  wire[27:0] T103;
  wire[31:0] T104;
  wire[31:0] T105;
  wire[31:0] T106;
  wire[23:0] T107;
  wire[31:0] T108;
  wire[31:0] T109;
  wire[31:0] T110;
  wire[15:0] T111;
  wire[31:0] T112;
  wire[31:0] T113;
  wire[31:0] T246;
  wire[15:0] T114;
  wire[31:0] T115;
  wire[31:0] T247;
  wire[23:0] T116;
  wire[31:0] T117;
  wire[31:0] T248;
  wire[27:0] T118;
  wire[31:0] T119;
  wire[31:0] T249;
  wire[29:0] T120;
  wire[31:0] T121;
  wire[31:0] T250;
  wire[30:0] T122;
  wire T123;
  wire T124;
  wire T125;
  wire T126;
  wire T127;
  wire T128;
  wire[55:0] adjustedSig;
  wire T129;
  wire[55:0] T130;
  wire[55:0] T131;
  wire[55:0] T132;
  wire common_totalUnderflow;
  wire T133;
  wire[15:0] T134;
  wire[14:0] T251;
  wire[3:0] T135;
  wire[3:0] T136;
  wire[2:0] T137;
  wire[55:0] T138;
  wire[54:0] T139;
  wire[54:0] T140;
  wire[54:0] T141;
  wire T142;
  wire roundingMode_odd;
  wire[54:0] T252;
  wire[53:0] T143;
  wire[55:0] T144;
  wire[55:0] T145;
  wire[55:0] T146;
  wire[54:0] T147;
  wire[54:0] T148;
  wire[54:0] T149;
  wire T150;
  wire T151;
  wire T152;
  wire roundingMode_near_even;
  wire[55:0] T153;
  wire[54:0] T253;
  wire[53:0] T154;
  wire[55:0] T155;
  wire T156;
  wire T157;
  wire roundMagUp;
  wire T158;
  wire T159;
  wire roundingMode_max;
  wire T160;
  wire roundingMode_min;
  wire T161;
  wire T162;
  wire roundingMode_near_maxMag;
  wire[10:0] T254;
  wire T255;
  wire[13:0] T256;
  wire T257;
  wire commonCase;
  wire T163;
  wire T164;
  wire T165;
  wire notNaN_isSpecialInfOut;
  wire T166;
  wire isNaNOut;
  wire underflow;
  wire common_underflow;
  wire T167;
  wire T168;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire T173;
  wire T174;
  wire[1:0] T175;
  wire T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  wire T182;
  wire T183;
  wire T184;
  wire T185;
  wire T186;
  wire T187;
  wire T188;
  wire T189;
  wire T190;
  wire T191;
  wire T192;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  wire T198;
  wire T199;
  wire[1:0] T200;
  wire overflow;
  wire common_overflow;
  wire T201;
  wire[5:0] T202;
  wire[1:0] T203;
  wire[64:0] T204;
  wire[63:0] T205;
  wire[51:0] fractOut;
  wire[51:0] T206;
  wire[51:0] T258;
  wire pegMaxFiniteMagOut;
  wire T207;
  wire overflow_roundMagUp;
  wire T208;
  wire[51:0] T209;
  wire[51:0] common_fractOut;
  wire[51:0] T210;
  wire[51:0] T211;
  wire[51:0] T212;
  wire[51:0] T213;
  wire T214;
  wire T215;
  wire[11:0] expOut;
  wire[11:0] T216;
  wire[11:0] T217;
  wire[11:0] T218;
  wire notNaN_isInfOut;
  wire T219;
  wire[11:0] T220;
  wire[11:0] T221;
  wire[11:0] T222;
  wire[11:0] T223;
  wire pegMinNonzeroMagOut;
  wire T224;
  wire T225;
  wire[11:0] T226;
  wire[11:0] T227;
  wire[11:0] T228;
  wire[11:0] T229;
  wire[11:0] T230;
  wire[11:0] T231;
  wire[11:0] T232;
  wire[11:0] T233;
  wire[11:0] T234;
  wire[11:0] T235;
  wire[11:0] T236;
  wire[11:0] T237;
  wire T238;
  wire[11:0] common_expOut;
  wire[11:0] T239;
  wire signOut;


  assign io_exceptionFlags = T0;
  assign T0 = {T203, T1};
  assign T1 = {overflow, T2};
  assign T2 = {underflow, inexact};
  assign inexact = overflow | T3;
  assign T3 = commonCase & common_inexact;
  assign common_inexact = T4;
  assign T4 = common_totalUnderflow | T5;
  assign T5 = T129 | T6;
  assign T6 = T7 != 56'h0;
  assign T7 = adjustedSig & T8;
  assign T8 = {1'h0, T9};
  assign T9 = T10 >> 1'h1;
  assign T10 = {T11, 2'h3};
  assign T11 = T12 | T240;
  assign T240 = {53'h0, doShiftSigDown1};
  assign doShiftSigDown1 = adjustedSig[55];
  assign T12 = T128 ? T13 : 54'h0;
  assign T13 = T127 ? T38 : T241;
  assign T241 = {51'h0, T14};
  assign T14 = T37 ? T15 : 3'h0;
  assign T15 = T36 ? T16 : 3'h0;
  assign T16 = T35 ? T17 : 3'h0;
  assign T17 = T34 ? T18 : 3'h0;
  assign T18 = {T30, T19};
  assign T19 = T20[2];
  assign T20 = T21[2:0];
  assign T21 = $signed(65'h10000000000000000) >>> T22;
  assign T22 = T23[5:0];
  assign T23 = T24[6:0];
  assign T24 = T25[7:0];
  assign T25 = T26[8:0];
  assign T26 = T27[9:0];
  assign T27 = T28[10:0];
  assign T28 = ~ T29;
  assign T29 = io_in_sExp[11:0];
  assign T30 = {T33, T31};
  assign T31 = T32[1];
  assign T32 = T20[1:0];
  assign T33 = T32[0];
  assign T34 = T23[6];
  assign T35 = T24[7];
  assign T36 = T25[8];
  assign T37 = T26[9];
  assign T38 = {T39, 3'h7};
  assign T39 = ~ T40;
  assign T40 = T126 ? 51'h0 : T41;
  assign T41 = ~ T42;
  assign T42 = ~ T43;
  assign T43 = T125 ? 51'h0 : T44;
  assign T44 = ~ T45;
  assign T45 = ~ T46;
  assign T46 = T124 ? 51'h0 : T47;
  assign T47 = ~ T48;
  assign T48 = ~ T49;
  assign T49 = T123 ? 51'h0 : T50;
  assign T50 = ~ T51;
  assign T51 = {T92, T52};
  assign T52 = {T67, T53};
  assign T53 = {T63, T54};
  assign T54 = T55[2];
  assign T55 = T56[18:16];
  assign T56 = T57[50:32];
  assign T57 = T58[63:13];
  assign T58 = $signed(65'h10000000000000000) >>> T59;
  assign T59 = T60[5:0];
  assign T60 = T61[6:0];
  assign T61 = T62[7:0];
  assign T62 = T26[8:0];
  assign T63 = {T66, T64};
  assign T64 = T65[1];
  assign T65 = T55[1:0];
  assign T66 = T65[0];
  assign T67 = T90 | T68;
  assign T68 = T69 & 16'haaaa;
  assign T69 = T70 << 1'h1;
  assign T70 = T71[14:0];
  assign T71 = T88 | T72;
  assign T72 = T73 & 16'hcccc;
  assign T73 = T74 << 2'h2;
  assign T74 = T75[13:0];
  assign T75 = T86 | T76;
  assign T76 = T77 & 16'hf0f0;
  assign T77 = T78 << 3'h4;
  assign T78 = T79[11:0];
  assign T79 = T84 | T80;
  assign T80 = T81 & 16'hff00;
  assign T81 = T82 << 4'h8;
  assign T82 = T83[7:0];
  assign T83 = T56[15:0];
  assign T84 = T242 & 16'hff;
  assign T242 = {8'h0, T85};
  assign T85 = T83 >> 4'h8;
  assign T86 = T243 & 16'hf0f;
  assign T243 = {4'h0, T87};
  assign T87 = T79 >> 3'h4;
  assign T88 = T244 & 16'h3333;
  assign T244 = {2'h0, T89};
  assign T89 = T75 >> 2'h2;
  assign T90 = T245 & 16'h5555;
  assign T245 = {1'h0, T91};
  assign T91 = T71 >> 1'h1;
  assign T92 = T121 | T93;
  assign T93 = T94 & 32'haaaaaaaa;
  assign T94 = T95 << 1'h1;
  assign T95 = T96[30:0];
  assign T96 = T119 | T97;
  assign T97 = T98 & 32'hcccccccc;
  assign T98 = T99 << 2'h2;
  assign T99 = T100[29:0];
  assign T100 = T117 | T101;
  assign T101 = T102 & 32'hf0f0f0f0;
  assign T102 = T103 << 3'h4;
  assign T103 = T104[27:0];
  assign T104 = T115 | T105;
  assign T105 = T106 & 32'hff00ff00;
  assign T106 = T107 << 4'h8;
  assign T107 = T108[23:0];
  assign T108 = T113 | T109;
  assign T109 = T110 & 32'hffff0000;
  assign T110 = T111 << 5'h10;
  assign T111 = T112[15:0];
  assign T112 = T57[31:0];
  assign T113 = T246 & 32'hffff;
  assign T246 = {16'h0, T114};
  assign T114 = T112 >> 5'h10;
  assign T115 = T247 & 32'hff00ff;
  assign T247 = {8'h0, T116};
  assign T116 = T108 >> 4'h8;
  assign T117 = T248 & 32'hf0f0f0f;
  assign T248 = {4'h0, T118};
  assign T118 = T104 >> 3'h4;
  assign T119 = T249 & 32'h33333333;
  assign T249 = {2'h0, T120};
  assign T120 = T100 >> 2'h2;
  assign T121 = T250 & 32'h55555555;
  assign T250 = {1'h0, T122};
  assign T122 = T96 >> 1'h1;
  assign T123 = T60[6];
  assign T124 = T61[7];
  assign T125 = T62[8];
  assign T126 = T26[9];
  assign T127 = T27[10];
  assign T128 = T28[11];
  assign adjustedSig = io_in_sig << 1'h0;
  assign T129 = T130 != 56'h0;
  assign T130 = adjustedSig & T131;
  assign T131 = T132 & T10;
  assign T132 = ~ T8;
  assign common_totalUnderflow = T133;
  assign T133 = $signed(T134) < $signed(11'h3ce);
  assign T134 = T256 + T251;
  assign T251 = {T254, T135};
  assign T135 = T136;
  assign T136 = {1'h0, T137};
  assign T137 = T138 >> 6'h35;
  assign T138 = T156 ? T146 : T139;
  assign T139 = T252 | T140;
  assign T140 = T142 ? T141 : 55'h0;
  assign T141 = T131 >> 1'h1;
  assign T142 = roundingMode_odd & T5;
  assign roundingMode_odd = io_roundingMode == 3'h6;
  assign T252 = {1'h0, T143};
  assign T143 = T144 >> 2'h2;
  assign T144 = adjustedSig & T145;
  assign T145 = ~ T10;
  assign T146 = T153 & T147;
  assign T147 = ~ T148;
  assign T148 = T150 ? T149 : 55'h0;
  assign T149 = T10 >> 1'h1;
  assign T150 = T152 & T151;
  assign T151 = T6 ^ 1'h1;
  assign T152 = roundingMode_near_even & T129;
  assign roundingMode_near_even = io_roundingMode == 3'h0;
  assign T153 = T253 + 55'h1;
  assign T253 = {1'h0, T154};
  assign T154 = T155 >> 2'h2;
  assign T155 = adjustedSig | T10;
  assign T156 = T161 | T157;
  assign T157 = roundMagUp & T5;
  assign roundMagUp = T160 | T158;
  assign T158 = roundingMode_max & T159;
  assign T159 = io_in_sign ^ 1'h1;
  assign roundingMode_max = io_roundingMode == 3'h3;
  assign T160 = roundingMode_min & io_in_sign;
  assign roundingMode_min = io_roundingMode == 3'h2;
  assign T161 = T162 & T129;
  assign T162 = roundingMode_near_even | roundingMode_near_maxMag;
  assign roundingMode_near_maxMag = io_roundingMode == 3'h4;
  assign T254 = T255 ? 11'h7ff : 11'h0;
  assign T255 = T135[2];
  assign T256 = {T257, io_in_sExp};
  assign T257 = io_in_sExp[12];
  assign commonCase = T164 & T163;
  assign T163 = io_in_isZero ^ 1'h1;
  assign T164 = T166 & T165;
  assign T165 = notNaN_isSpecialInfOut ^ 1'h1;
  assign notNaN_isSpecialInfOut = io_infiniteExc | io_in_isInf;
  assign T166 = isNaNOut ^ 1'h1;
  assign isNaNOut = io_invalidExc | io_in_isNaN;
  assign underflow = commonCase & common_underflow;
  assign common_underflow = T167;
  assign T167 = common_totalUnderflow | T168;
  assign T168 = T194 & T169;
  assign T169 = T170 ^ 1'h1;
  assign T170 = T183 & T171;
  assign T171 = T178 | T172;
  assign T172 = roundMagUp & T173;
  assign T173 = T176 | T174;
  assign T174 = T175 != 2'h0;
  assign T175 = adjustedSig[1:0];
  assign T176 = doShiftSigDown1 & T177;
  assign T177 = adjustedSig[2];
  assign T178 = T182 & T179;
  assign T179 = doShiftSigDown1 ? T181 : T180;
  assign T180 = adjustedSig[1];
  assign T181 = adjustedSig[2];
  assign T182 = roundingMode_near_even | roundingMode_near_maxMag;
  assign T183 = T184 & T129;
  assign T184 = T188 & T185;
  assign T185 = doShiftSigDown1 ? T187 : T186;
  assign T186 = T138[53];
  assign T187 = T138[54];
  assign T188 = T193 & T189;
  assign T189 = T190 ^ 1'h1;
  assign T190 = doShiftSigDown1 ? T192 : T191;
  assign T191 = T10[3];
  assign T192 = T10[4];
  assign T193 = io_detectTininess == 1'h1;
  assign T194 = T198 & T195;
  assign T195 = doShiftSigDown1 ? T197 : T196;
  assign T196 = T10[2];
  assign T197 = T10[3];
  assign T198 = T5 & T199;
  assign T199 = $signed(T200) <= $signed(1'h0);
  assign T200 = $signed(io_in_sExp) >>> 4'hb;
  assign overflow = commonCase & common_overflow;
  assign common_overflow = T201;
  assign T201 = $signed(3'h3) <= $signed(T202);
  assign T202 = $signed(T134) >>> 4'ha;
  assign T203 = {io_invalidExc, io_infiniteExc};
  assign io_out = T204;
  assign T204 = {signOut, T205};
  assign T205 = {expOut, fractOut};
  assign fractOut = T209 | T206;
  assign T206 = 52'h0 - T258;
  assign T258 = {51'h0, pegMaxFiniteMagOut};
  assign pegMaxFiniteMagOut = overflow & T207;
  assign T207 = overflow_roundMagUp ^ 1'h1;
  assign overflow_roundMagUp = T208 | roundMagUp;
  assign T208 = roundingMode_near_even | roundingMode_near_maxMag;
  assign T209 = T214 ? T213 : common_fractOut;
  assign common_fractOut = T210;
  assign T210 = doShiftSigDown1 ? T212 : T211;
  assign T211 = T138[51:0];
  assign T212 = T138[52:1];
  assign T213 = isNaNOut ? 52'h8000000000000 : 52'h0;
  assign T214 = T215 | common_totalUnderflow;
  assign T215 = isNaNOut | io_in_isZero;
  assign expOut = T217 | T216;
  assign T216 = isNaNOut ? 12'he00 : 12'h0;
  assign T217 = T220 | T218;
  assign T218 = notNaN_isInfOut ? 12'hc00 : 12'h0;
  assign notNaN_isInfOut = notNaN_isSpecialInfOut | T219;
  assign T219 = overflow & overflow_roundMagUp;
  assign T220 = T222 | T221;
  assign T221 = pegMaxFiniteMagOut ? 12'hbff : 12'h0;
  assign T222 = T226 | T223;
  assign T223 = pegMinNonzeroMagOut ? 12'h3ce : 12'h0;
  assign pegMinNonzeroMagOut = T225 & T224;
  assign T224 = roundMagUp | roundingMode_odd;
  assign T225 = commonCase & common_totalUnderflow;
  assign T226 = T229 & T227;
  assign T227 = ~ T228;
  assign T228 = notNaN_isInfOut ? 12'h200 : 12'h0;
  assign T229 = T232 & T230;
  assign T230 = ~ T231;
  assign T231 = pegMaxFiniteMagOut ? 12'h400 : 12'h0;
  assign T232 = T235 & T233;
  assign T233 = ~ T234;
  assign T234 = pegMinNonzeroMagOut ? 12'hc31 : 12'h0;
  assign T235 = common_expOut & T236;
  assign T236 = ~ T237;
  assign T237 = T238 ? 12'he00 : 12'h0;
  assign T238 = io_in_isZero | common_totalUnderflow;
  assign common_expOut = T239;
  assign T239 = T134[11:0];
  assign signOut = isNaNOut ? 1'h0 : io_in_sign;
endmodule

module RoundRawFNToRecFN(
    input  io_invalidExc,
    input  io_infiniteExc,
    input  io_in_isNaN,
    input  io_in_isInf,
    input  io_in_isZero,
    input  io_in_sign,
    input [12:0] io_in_sExp,
    input [55:0] io_in_sig,
    input [2:0] io_roundingMode,
    input  io_detectTininess,
    output[64:0] io_out,
    output[4:0] io_exceptionFlags
);

  wire[64:0] roundAnyRawFNToRecFN_io_out;
  wire[4:0] roundAnyRawFNToRecFN_io_exceptionFlags;


  assign io_exceptionFlags = roundAnyRawFNToRecFN_io_exceptionFlags;
  assign io_out = roundAnyRawFNToRecFN_io_out;
  RoundAnyRawFNToRecFN roundAnyRawFNToRecFN(
       .io_invalidExc( io_invalidExc ),
       .io_infiniteExc( io_infiniteExc ),
       .io_in_isNaN( io_in_isNaN ),
       .io_in_isInf( io_in_isInf ),
       .io_in_isZero( io_in_isZero ),
       .io_in_sign( io_in_sign ),
       .io_in_sExp( io_in_sExp ),
       .io_in_sig( io_in_sig ),
       .io_roundingMode( io_roundingMode ),
       .io_detectTininess( io_detectTininess ),
       .io_out( roundAnyRawFNToRecFN_io_out ),
       .io_exceptionFlags( roundAnyRawFNToRecFN_io_exceptionFlags )
  );
endmodule

module MulAddRecFN(
    input [1:0] io_op,
    input [64:0] io_a,
    input [64:0] io_b,
    input [64:0] io_c,
    input [2:0] io_roundingMode,
    input  io_detectTininess,
    output[64:0] io_out,
    output[4:0] io_exceptionFlags
);

  wire[106:0] mulAddResult;
  wire[106:0] T1;
  wire[106:0] T2;
  wire[105:0] T0;
  wire[52:0] mulAddRecFNToRaw_preMul_io_mulAddA;
  wire[52:0] mulAddRecFNToRaw_preMul_io_mulAddB;
  wire[105:0] mulAddRecFNToRaw_preMul_io_mulAddC;
  wire mulAddRecFNToRaw_preMul_io_toPostMul_isSigNaNAny;
  wire mulAddRecFNToRaw_preMul_io_toPostMul_isNaNAOrB;
  wire mulAddRecFNToRaw_preMul_io_toPostMul_isInfA;
  wire mulAddRecFNToRaw_preMul_io_toPostMul_isZeroA;
  wire mulAddRecFNToRaw_preMul_io_toPostMul_isInfB;
  wire mulAddRecFNToRaw_preMul_io_toPostMul_isZeroB;
  wire mulAddRecFNToRaw_preMul_io_toPostMul_signProd;
  wire mulAddRecFNToRaw_preMul_io_toPostMul_isNaNC;
  wire mulAddRecFNToRaw_preMul_io_toPostMul_isInfC;
  wire mulAddRecFNToRaw_preMul_io_toPostMul_isZeroC;
  wire[12:0] mulAddRecFNToRaw_preMul_io_toPostMul_sExpSum;
  wire mulAddRecFNToRaw_preMul_io_toPostMul_doSubMags;
  wire mulAddRecFNToRaw_preMul_io_toPostMul_CIsDominant;
  wire[5:0] mulAddRecFNToRaw_preMul_io_toPostMul_CDom_CAlignDist;
  wire[54:0] mulAddRecFNToRaw_preMul_io_toPostMul_highAlignedSigC;
  wire mulAddRecFNToRaw_preMul_io_toPostMul_bit0AlignedSigC;
  wire mulAddRecFNToRaw_postMul_io_invalidExc;
  wire mulAddRecFNToRaw_postMul_io_rawOut_isNaN;
  wire mulAddRecFNToRaw_postMul_io_rawOut_isInf;
  wire mulAddRecFNToRaw_postMul_io_rawOut_isZero;
  wire mulAddRecFNToRaw_postMul_io_rawOut_sign;
  wire[12:0] mulAddRecFNToRaw_postMul_io_rawOut_sExp;
  wire[55:0] mulAddRecFNToRaw_postMul_io_rawOut_sig;
  wire[64:0] roundRawFNToRecFN_io_out;
  wire[4:0] roundRawFNToRecFN_io_exceptionFlags;


  assign mulAddResult = T2 + T1;
  assign T1 = {1'h0, mulAddRecFNToRaw_preMul_io_mulAddC};
  assign T2 = {1'h0, T0};
  assign T0 = mulAddRecFNToRaw_preMul_io_mulAddA * mulAddRecFNToRaw_preMul_io_mulAddB;
  assign io_exceptionFlags = roundRawFNToRecFN_io_exceptionFlags;
  assign io_out = roundRawFNToRecFN_io_out;
  MulAddRecFNToRaw_preMul mulAddRecFNToRaw_preMul(
       .io_op( io_op ),
       .io_a( io_a ),
       .io_b( io_b ),
       .io_c( io_c ),
       .io_mulAddA( mulAddRecFNToRaw_preMul_io_mulAddA ),
       .io_mulAddB( mulAddRecFNToRaw_preMul_io_mulAddB ),
       .io_mulAddC( mulAddRecFNToRaw_preMul_io_mulAddC ),
       .io_toPostMul_isSigNaNAny( mulAddRecFNToRaw_preMul_io_toPostMul_isSigNaNAny ),
       .io_toPostMul_isNaNAOrB( mulAddRecFNToRaw_preMul_io_toPostMul_isNaNAOrB ),
       .io_toPostMul_isInfA( mulAddRecFNToRaw_preMul_io_toPostMul_isInfA ),
       .io_toPostMul_isZeroA( mulAddRecFNToRaw_preMul_io_toPostMul_isZeroA ),
       .io_toPostMul_isInfB( mulAddRecFNToRaw_preMul_io_toPostMul_isInfB ),
       .io_toPostMul_isZeroB( mulAddRecFNToRaw_preMul_io_toPostMul_isZeroB ),
       .io_toPostMul_signProd( mulAddRecFNToRaw_preMul_io_toPostMul_signProd ),
       .io_toPostMul_isNaNC( mulAddRecFNToRaw_preMul_io_toPostMul_isNaNC ),
       .io_toPostMul_isInfC( mulAddRecFNToRaw_preMul_io_toPostMul_isInfC ),
       .io_toPostMul_isZeroC( mulAddRecFNToRaw_preMul_io_toPostMul_isZeroC ),
       .io_toPostMul_sExpSum( mulAddRecFNToRaw_preMul_io_toPostMul_sExpSum ),
       .io_toPostMul_doSubMags( mulAddRecFNToRaw_preMul_io_toPostMul_doSubMags ),
       .io_toPostMul_CIsDominant( mulAddRecFNToRaw_preMul_io_toPostMul_CIsDominant ),
       .io_toPostMul_CDom_CAlignDist( mulAddRecFNToRaw_preMul_io_toPostMul_CDom_CAlignDist ),
       .io_toPostMul_highAlignedSigC( mulAddRecFNToRaw_preMul_io_toPostMul_highAlignedSigC ),
       .io_toPostMul_bit0AlignedSigC( mulAddRecFNToRaw_preMul_io_toPostMul_bit0AlignedSigC )
  );
  MulAddRecFNToRaw_postMul mulAddRecFNToRaw_postMul(
       .io_fromPreMul_isSigNaNAny( mulAddRecFNToRaw_preMul_io_toPostMul_isSigNaNAny ),
       .io_fromPreMul_isNaNAOrB( mulAddRecFNToRaw_preMul_io_toPostMul_isNaNAOrB ),
       .io_fromPreMul_isInfA( mulAddRecFNToRaw_preMul_io_toPostMul_isInfA ),
       .io_fromPreMul_isZeroA( mulAddRecFNToRaw_preMul_io_toPostMul_isZeroA ),
       .io_fromPreMul_isInfB( mulAddRecFNToRaw_preMul_io_toPostMul_isInfB ),
       .io_fromPreMul_isZeroB( mulAddRecFNToRaw_preMul_io_toPostMul_isZeroB ),
       .io_fromPreMul_signProd( mulAddRecFNToRaw_preMul_io_toPostMul_signProd ),
       .io_fromPreMul_isNaNC( mulAddRecFNToRaw_preMul_io_toPostMul_isNaNC ),
       .io_fromPreMul_isInfC( mulAddRecFNToRaw_preMul_io_toPostMul_isInfC ),
       .io_fromPreMul_isZeroC( mulAddRecFNToRaw_preMul_io_toPostMul_isZeroC ),
       .io_fromPreMul_sExpSum( mulAddRecFNToRaw_preMul_io_toPostMul_sExpSum ),
       .io_fromPreMul_doSubMags( mulAddRecFNToRaw_preMul_io_toPostMul_doSubMags ),
       .io_fromPreMul_CIsDominant( mulAddRecFNToRaw_preMul_io_toPostMul_CIsDominant ),
       .io_fromPreMul_CDom_CAlignDist( mulAddRecFNToRaw_preMul_io_toPostMul_CDom_CAlignDist ),
       .io_fromPreMul_highAlignedSigC( mulAddRecFNToRaw_preMul_io_toPostMul_highAlignedSigC ),
       .io_fromPreMul_bit0AlignedSigC( mulAddRecFNToRaw_preMul_io_toPostMul_bit0AlignedSigC ),
       .io_mulAddResult( mulAddResult ),
       .io_roundingMode( io_roundingMode ),
       .io_invalidExc( mulAddRecFNToRaw_postMul_io_invalidExc ),
       .io_rawOut_isNaN( mulAddRecFNToRaw_postMul_io_rawOut_isNaN ),
       .io_rawOut_isInf( mulAddRecFNToRaw_postMul_io_rawOut_isInf ),
       .io_rawOut_isZero( mulAddRecFNToRaw_postMul_io_rawOut_isZero ),
       .io_rawOut_sign( mulAddRecFNToRaw_postMul_io_rawOut_sign ),
       .io_rawOut_sExp( mulAddRecFNToRaw_postMul_io_rawOut_sExp ),
       .io_rawOut_sig( mulAddRecFNToRaw_postMul_io_rawOut_sig )
  );
  RoundRawFNToRecFN roundRawFNToRecFN(
       .io_invalidExc( mulAddRecFNToRaw_postMul_io_invalidExc ),
       .io_infiniteExc( 1'h0 ),
       .io_in_isNaN( mulAddRecFNToRaw_postMul_io_rawOut_isNaN ),
       .io_in_isInf( mulAddRecFNToRaw_postMul_io_rawOut_isInf ),
       .io_in_isZero( mulAddRecFNToRaw_postMul_io_rawOut_isZero ),
       .io_in_sign( mulAddRecFNToRaw_postMul_io_rawOut_sign ),
       .io_in_sExp( mulAddRecFNToRaw_postMul_io_rawOut_sExp ),
       .io_in_sig( mulAddRecFNToRaw_postMul_io_rawOut_sig ),
       .io_roundingMode( io_roundingMode ),
       .io_detectTininess( io_detectTininess ),
       .io_out( roundRawFNToRecFN_io_out ),
       .io_exceptionFlags( roundRawFNToRecFN_io_exceptionFlags )
  );
endmodule

module ValExec_MulAddRecF64_add(
    input [63:0] io_a,
    input [63:0] io_b,
    input [2:0] io_roundingMode,
    input  io_detectTininess,
    input [63:0] io_expected_out,
    input [4:0] io_expected_exceptionFlags,
    output[64:0] io_expected_recOut,
    output[64:0] io_actual_out,
    output[4:0] io_actual_exceptionFlags,
    output io_check,
    output io_pass
);

  wire[64:0] T0;
  wire[60:0] T1;
  wire[51:0] T2;
  wire[53:0] T3;
  wire[53:0] T4;
  wire[52:0] T5;
  wire[51:0] T6;
  wire[51:0] T7;
  wire[51:0] T8;
  wire[50:0] T9;
  wire[114:0] T10;
  wire[5:0] T344;
  wire[5:0] T345;
  wire[5:0] T346;
  wire[5:0] T347;
  wire[5:0] T348;
  wire[5:0] T349;
  wire[5:0] T350;
  wire[5:0] T351;
  wire[5:0] T352;
  wire[5:0] T353;
  wire[5:0] T354;
  wire[5:0] T355;
  wire[5:0] T356;
  wire[5:0] T357;
  wire[5:0] T358;
  wire[5:0] T359;
  wire[5:0] T360;
  wire[5:0] T361;
  wire[5:0] T362;
  wire[5:0] T363;
  wire[5:0] T364;
  wire[5:0] T365;
  wire[5:0] T366;
  wire[5:0] T367;
  wire[5:0] T368;
  wire[5:0] T369;
  wire[5:0] T370;
  wire[5:0] T371;
  wire[5:0] T372;
  wire[5:0] T373;
  wire[5:0] T374;
  wire[5:0] T375;
  wire[5:0] T376;
  wire[5:0] T377;
  wire[5:0] T378;
  wire[5:0] T379;
  wire[5:0] T380;
  wire[5:0] T381;
  wire[5:0] T382;
  wire[5:0] T383;
  wire[5:0] T384;
  wire[5:0] T385;
  wire[5:0] T386;
  wire[5:0] T387;
  wire[5:0] T388;
  wire[5:0] T389;
  wire[5:0] T390;
  wire[5:0] T391;
  wire[5:0] T392;
  wire[5:0] T393;
  wire[5:0] T394;
  wire T395;
  wire[51:0] T12;
  wire[19:0] T13;
  wire[3:0] T14;
  wire[1:0] T15;
  wire T16;
  wire[1:0] T17;
  wire[3:0] T18;
  wire[19:0] T19;
  wire T20;
  wire[1:0] T21;
  wire T22;
  wire[1:0] T23;
  wire T24;
  wire[15:0] T25;
  wire[15:0] T26;
  wire[15:0] T27;
  wire[14:0] T28;
  wire[15:0] T29;
  wire[15:0] T30;
  wire[15:0] T31;
  wire[13:0] T32;
  wire[15:0] T33;
  wire[15:0] T34;
  wire[15:0] T35;
  wire[11:0] T36;
  wire[15:0] T37;
  wire[15:0] T38;
  wire[15:0] T39;
  wire[7:0] T40;
  wire[15:0] T41;
  wire[15:0] T42;
  wire[15:0] T396;
  wire[7:0] T43;
  wire[15:0] T44;
  wire[15:0] T397;
  wire[11:0] T45;
  wire[15:0] T46;
  wire[15:0] T398;
  wire[13:0] T47;
  wire[15:0] T48;
  wire[15:0] T399;
  wire[14:0] T49;
  wire[31:0] T50;
  wire[31:0] T51;
  wire[31:0] T52;
  wire[30:0] T53;
  wire[31:0] T54;
  wire[31:0] T55;
  wire[31:0] T56;
  wire[29:0] T57;
  wire[31:0] T58;
  wire[31:0] T59;
  wire[31:0] T60;
  wire[27:0] T61;
  wire[31:0] T62;
  wire[31:0] T63;
  wire[31:0] T64;
  wire[23:0] T65;
  wire[31:0] T66;
  wire[31:0] T67;
  wire[31:0] T68;
  wire[15:0] T69;
  wire[31:0] T70;
  wire[31:0] T71;
  wire[31:0] T400;
  wire[15:0] T72;
  wire[31:0] T73;
  wire[31:0] T401;
  wire[23:0] T74;
  wire[31:0] T75;
  wire[31:0] T402;
  wire[27:0] T76;
  wire[31:0] T77;
  wire[31:0] T403;
  wire[29:0] T78;
  wire[31:0] T79;
  wire[31:0] T404;
  wire[30:0] T80;
  wire T405;
  wire T406;
  wire T407;
  wire T408;
  wire T409;
  wire T410;
  wire T411;
  wire T412;
  wire T413;
  wire T414;
  wire T415;
  wire T416;
  wire T417;
  wire T418;
  wire T419;
  wire T420;
  wire T421;
  wire T422;
  wire T423;
  wire T424;
  wire T425;
  wire T426;
  wire T427;
  wire T428;
  wire T429;
  wire T430;
  wire T431;
  wire T432;
  wire T433;
  wire T434;
  wire T435;
  wire T436;
  wire T437;
  wire T438;
  wire T439;
  wire T440;
  wire T441;
  wire T442;
  wire T443;
  wire T444;
  wire T445;
  wire T446;
  wire T447;
  wire T448;
  wire T449;
  wire T450;
  wire T451;
  wire T452;
  wire T453;
  wire T454;
  wire T81;
  wire[10:0] T82;
  wire T83;
  wire T84;
  wire T85;
  wire[8:0] T86;
  wire[12:0] T87;
  wire[12:0] T88;
  wire[12:0] T89;
  wire[11:0] T90;
  wire[11:0] T91;
  wire[11:0] T455;
  wire[10:0] T92;
  wire[10:0] T456;
  wire[1:0] T93;
  wire[11:0] T94;
  wire[11:0] T457;
  wire[11:0] T95;
  wire[11:0] T458;
  wire[3:0] T96;
  wire[2:0] T97;
  wire[2:0] T459;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire[1:0] T102;
  wire[2:0] T103;
  wire[2:0] T104;
  wire T105;
  wire T106;
  wire T107;
  wire[64:0] T108;
  wire[60:0] T109;
  wire[51:0] T110;
  wire[53:0] T111;
  wire[53:0] T112;
  wire[52:0] T113;
  wire[51:0] T114;
  wire[51:0] T115;
  wire[51:0] T116;
  wire[50:0] T117;
  wire[114:0] T118;
  wire[5:0] T460;
  wire[5:0] T461;
  wire[5:0] T462;
  wire[5:0] T463;
  wire[5:0] T464;
  wire[5:0] T465;
  wire[5:0] T466;
  wire[5:0] T467;
  wire[5:0] T468;
  wire[5:0] T469;
  wire[5:0] T470;
  wire[5:0] T471;
  wire[5:0] T472;
  wire[5:0] T473;
  wire[5:0] T474;
  wire[5:0] T475;
  wire[5:0] T476;
  wire[5:0] T477;
  wire[5:0] T478;
  wire[5:0] T479;
  wire[5:0] T480;
  wire[5:0] T481;
  wire[5:0] T482;
  wire[5:0] T483;
  wire[5:0] T484;
  wire[5:0] T485;
  wire[5:0] T486;
  wire[5:0] T487;
  wire[5:0] T488;
  wire[5:0] T489;
  wire[5:0] T490;
  wire[5:0] T491;
  wire[5:0] T492;
  wire[5:0] T493;
  wire[5:0] T494;
  wire[5:0] T495;
  wire[5:0] T496;
  wire[5:0] T497;
  wire[5:0] T498;
  wire[5:0] T499;
  wire[5:0] T500;
  wire[5:0] T501;
  wire[5:0] T502;
  wire[5:0] T503;
  wire[5:0] T504;
  wire[5:0] T505;
  wire[5:0] T506;
  wire[5:0] T507;
  wire[5:0] T508;
  wire[5:0] T509;
  wire[5:0] T510;
  wire T511;
  wire[51:0] T120;
  wire[19:0] T121;
  wire[3:0] T122;
  wire[1:0] T123;
  wire T124;
  wire[1:0] T125;
  wire[3:0] T126;
  wire[19:0] T127;
  wire T128;
  wire[1:0] T129;
  wire T130;
  wire[1:0] T131;
  wire T132;
  wire[15:0] T133;
  wire[15:0] T134;
  wire[15:0] T135;
  wire[14:0] T136;
  wire[15:0] T137;
  wire[15:0] T138;
  wire[15:0] T139;
  wire[13:0] T140;
  wire[15:0] T141;
  wire[15:0] T142;
  wire[15:0] T143;
  wire[11:0] T144;
  wire[15:0] T145;
  wire[15:0] T146;
  wire[15:0] T147;
  wire[7:0] T148;
  wire[15:0] T149;
  wire[15:0] T150;
  wire[15:0] T512;
  wire[7:0] T151;
  wire[15:0] T152;
  wire[15:0] T513;
  wire[11:0] T153;
  wire[15:0] T154;
  wire[15:0] T514;
  wire[13:0] T155;
  wire[15:0] T156;
  wire[15:0] T515;
  wire[14:0] T157;
  wire[31:0] T158;
  wire[31:0] T159;
  wire[31:0] T160;
  wire[30:0] T161;
  wire[31:0] T162;
  wire[31:0] T163;
  wire[31:0] T164;
  wire[29:0] T165;
  wire[31:0] T166;
  wire[31:0] T167;
  wire[31:0] T168;
  wire[27:0] T169;
  wire[31:0] T170;
  wire[31:0] T171;
  wire[31:0] T172;
  wire[23:0] T173;
  wire[31:0] T174;
  wire[31:0] T175;
  wire[31:0] T176;
  wire[15:0] T177;
  wire[31:0] T178;
  wire[31:0] T179;
  wire[31:0] T516;
  wire[15:0] T180;
  wire[31:0] T181;
  wire[31:0] T517;
  wire[23:0] T182;
  wire[31:0] T183;
  wire[31:0] T518;
  wire[27:0] T184;
  wire[31:0] T185;
  wire[31:0] T519;
  wire[29:0] T186;
  wire[31:0] T187;
  wire[31:0] T520;
  wire[30:0] T188;
  wire T521;
  wire T522;
  wire T523;
  wire T524;
  wire T525;
  wire T526;
  wire T527;
  wire T528;
  wire T529;
  wire T530;
  wire T531;
  wire T532;
  wire T533;
  wire T534;
  wire T535;
  wire T536;
  wire T537;
  wire T538;
  wire T539;
  wire T540;
  wire T541;
  wire T542;
  wire T543;
  wire T544;
  wire T545;
  wire T546;
  wire T547;
  wire T548;
  wire T549;
  wire T550;
  wire T551;
  wire T552;
  wire T553;
  wire T554;
  wire T555;
  wire T556;
  wire T557;
  wire T558;
  wire T559;
  wire T560;
  wire T561;
  wire T562;
  wire T563;
  wire T564;
  wire T565;
  wire T566;
  wire T567;
  wire T568;
  wire T569;
  wire T570;
  wire T189;
  wire[10:0] T190;
  wire T191;
  wire T192;
  wire T193;
  wire[8:0] T194;
  wire[12:0] T195;
  wire[12:0] T196;
  wire[12:0] T197;
  wire[11:0] T198;
  wire[11:0] T199;
  wire[11:0] T571;
  wire[10:0] T200;
  wire[10:0] T572;
  wire[1:0] T201;
  wire[11:0] T202;
  wire[11:0] T573;
  wire[11:0] T203;
  wire[11:0] T574;
  wire[3:0] T204;
  wire[2:0] T205;
  wire[2:0] T575;
  wire T206;
  wire T207;
  wire T208;
  wire T209;
  wire[1:0] T210;
  wire[2:0] T211;
  wire[2:0] T212;
  wire T213;
  wire T214;
  wire T215;
  wire T216;
  wire T217;
  wire T218;
  wire T219;
  wire T220;
  wire T221;
  wire[3:0] T222;
  wire[3:0] T223;
  wire T224;
  wire[2:0] T225;
  wire T226;
  wire T227;
  wire[51:0] T228;
  wire[51:0] T229;
  wire T230;
  wire T231;
  wire T232;
  wire[2:0] T233;
  wire T234;
  wire[2:0] T235;
  wire[64:0] T236;
  wire[60:0] T237;
  wire[51:0] T238;
  wire[53:0] T239;
  wire[53:0] T240;
  wire[52:0] T241;
  wire[51:0] T242;
  wire[51:0] T243;
  wire[51:0] T244;
  wire[50:0] T245;
  wire[114:0] T246;
  wire[5:0] T576;
  wire[5:0] T577;
  wire[5:0] T578;
  wire[5:0] T579;
  wire[5:0] T580;
  wire[5:0] T581;
  wire[5:0] T582;
  wire[5:0] T583;
  wire[5:0] T584;
  wire[5:0] T585;
  wire[5:0] T586;
  wire[5:0] T587;
  wire[5:0] T588;
  wire[5:0] T589;
  wire[5:0] T590;
  wire[5:0] T591;
  wire[5:0] T592;
  wire[5:0] T593;
  wire[5:0] T594;
  wire[5:0] T595;
  wire[5:0] T596;
  wire[5:0] T597;
  wire[5:0] T598;
  wire[5:0] T599;
  wire[5:0] T600;
  wire[5:0] T601;
  wire[5:0] T602;
  wire[5:0] T603;
  wire[5:0] T604;
  wire[5:0] T605;
  wire[5:0] T606;
  wire[5:0] T607;
  wire[5:0] T608;
  wire[5:0] T609;
  wire[5:0] T610;
  wire[5:0] T611;
  wire[5:0] T612;
  wire[5:0] T613;
  wire[5:0] T614;
  wire[5:0] T615;
  wire[5:0] T616;
  wire[5:0] T617;
  wire[5:0] T618;
  wire[5:0] T619;
  wire[5:0] T620;
  wire[5:0] T621;
  wire[5:0] T622;
  wire[5:0] T623;
  wire[5:0] T624;
  wire[5:0] T625;
  wire[5:0] T626;
  wire T627;
  wire[51:0] T248;
  wire[19:0] T249;
  wire[3:0] T250;
  wire[1:0] T251;
  wire T252;
  wire[1:0] T253;
  wire[3:0] T254;
  wire[19:0] T255;
  wire T256;
  wire[1:0] T257;
  wire T258;
  wire[1:0] T259;
  wire T260;
  wire[15:0] T261;
  wire[15:0] T262;
  wire[15:0] T263;
  wire[14:0] T264;
  wire[15:0] T265;
  wire[15:0] T266;
  wire[15:0] T267;
  wire[13:0] T268;
  wire[15:0] T269;
  wire[15:0] T270;
  wire[15:0] T271;
  wire[11:0] T272;
  wire[15:0] T273;
  wire[15:0] T274;
  wire[15:0] T275;
  wire[7:0] T276;
  wire[15:0] T277;
  wire[15:0] T278;
  wire[15:0] T628;
  wire[7:0] T279;
  wire[15:0] T280;
  wire[15:0] T629;
  wire[11:0] T281;
  wire[15:0] T282;
  wire[15:0] T630;
  wire[13:0] T283;
  wire[15:0] T284;
  wire[15:0] T631;
  wire[14:0] T285;
  wire[31:0] T286;
  wire[31:0] T287;
  wire[31:0] T288;
  wire[30:0] T289;
  wire[31:0] T290;
  wire[31:0] T291;
  wire[31:0] T292;
  wire[29:0] T293;
  wire[31:0] T294;
  wire[31:0] T295;
  wire[31:0] T296;
  wire[27:0] T297;
  wire[31:0] T298;
  wire[31:0] T299;
  wire[31:0] T300;
  wire[23:0] T301;
  wire[31:0] T302;
  wire[31:0] T303;
  wire[31:0] T304;
  wire[15:0] T305;
  wire[31:0] T306;
  wire[31:0] T307;
  wire[31:0] T632;
  wire[15:0] T308;
  wire[31:0] T309;
  wire[31:0] T633;
  wire[23:0] T310;
  wire[31:0] T311;
  wire[31:0] T634;
  wire[27:0] T312;
  wire[31:0] T313;
  wire[31:0] T635;
  wire[29:0] T314;
  wire[31:0] T315;
  wire[31:0] T636;
  wire[30:0] T316;
  wire T637;
  wire T638;
  wire T639;
  wire T640;
  wire T641;
  wire T642;
  wire T643;
  wire T644;
  wire T645;
  wire T646;
  wire T647;
  wire T648;
  wire T649;
  wire T650;
  wire T651;
  wire T652;
  wire T653;
  wire T654;
  wire T655;
  wire T656;
  wire T657;
  wire T658;
  wire T659;
  wire T660;
  wire T661;
  wire T662;
  wire T663;
  wire T664;
  wire T665;
  wire T666;
  wire T667;
  wire T668;
  wire T669;
  wire T670;
  wire T671;
  wire T672;
  wire T673;
  wire T674;
  wire T675;
  wire T676;
  wire T677;
  wire T678;
  wire T679;
  wire T680;
  wire T681;
  wire T682;
  wire T683;
  wire T684;
  wire T685;
  wire T686;
  wire T317;
  wire[10:0] T318;
  wire T319;
  wire T320;
  wire T321;
  wire[8:0] T322;
  wire[12:0] T323;
  wire[12:0] T324;
  wire[12:0] T325;
  wire[11:0] T326;
  wire[11:0] T327;
  wire[11:0] T687;
  wire[10:0] T328;
  wire[10:0] T688;
  wire[1:0] T329;
  wire[11:0] T330;
  wire[11:0] T689;
  wire[11:0] T331;
  wire[11:0] T690;
  wire[3:0] T332;
  wire[2:0] T333;
  wire[2:0] T691;
  wire T334;
  wire T335;
  wire T336;
  wire T337;
  wire[1:0] T338;
  wire[2:0] T339;
  wire[2:0] T340;
  wire T341;
  wire T342;
  wire T343;
  wire[64:0] mulAddRecFN_io_out;
  wire[4:0] mulAddRecFN_io_exceptionFlags;


  assign T0 = {T96, T1};
  assign T1 = {T86, T2};
  assign T2 = T3[51:0];
  assign T3 = T4;
  assign T4 = {1'h0, T5};
  assign T5 = {T83, T6};
  assign T6 = T81 ? T8 : T7;
  assign T7 = io_b[51:0];
  assign T8 = T9 << 1'h1;
  assign T9 = T10[50:0];
  assign T10 = T7 << T344;
  assign T344 = T454 ? 1'h0 : T345;
  assign T345 = T453 ? 1'h1 : T346;
  assign T346 = T452 ? 2'h2 : T347;
  assign T347 = T451 ? 2'h3 : T348;
  assign T348 = T450 ? 3'h4 : T349;
  assign T349 = T449 ? 3'h5 : T350;
  assign T350 = T448 ? 3'h6 : T351;
  assign T351 = T447 ? 3'h7 : T352;
  assign T352 = T446 ? 4'h8 : T353;
  assign T353 = T445 ? 4'h9 : T354;
  assign T354 = T444 ? 4'ha : T355;
  assign T355 = T443 ? 4'hb : T356;
  assign T356 = T442 ? 4'hc : T357;
  assign T357 = T441 ? 4'hd : T358;
  assign T358 = T440 ? 4'he : T359;
  assign T359 = T439 ? 4'hf : T360;
  assign T360 = T438 ? 5'h10 : T361;
  assign T361 = T437 ? 5'h11 : T362;
  assign T362 = T436 ? 5'h12 : T363;
  assign T363 = T435 ? 5'h13 : T364;
  assign T364 = T434 ? 5'h14 : T365;
  assign T365 = T433 ? 5'h15 : T366;
  assign T366 = T432 ? 5'h16 : T367;
  assign T367 = T431 ? 5'h17 : T368;
  assign T368 = T430 ? 5'h18 : T369;
  assign T369 = T429 ? 5'h19 : T370;
  assign T370 = T428 ? 5'h1a : T371;
  assign T371 = T427 ? 5'h1b : T372;
  assign T372 = T426 ? 5'h1c : T373;
  assign T373 = T425 ? 5'h1d : T374;
  assign T374 = T424 ? 5'h1e : T375;
  assign T375 = T423 ? 5'h1f : T376;
  assign T376 = T422 ? 6'h20 : T377;
  assign T377 = T421 ? 6'h21 : T378;
  assign T378 = T420 ? 6'h22 : T379;
  assign T379 = T419 ? 6'h23 : T380;
  assign T380 = T418 ? 6'h24 : T381;
  assign T381 = T417 ? 6'h25 : T382;
  assign T382 = T416 ? 6'h26 : T383;
  assign T383 = T415 ? 6'h27 : T384;
  assign T384 = T414 ? 6'h28 : T385;
  assign T385 = T413 ? 6'h29 : T386;
  assign T386 = T412 ? 6'h2a : T387;
  assign T387 = T411 ? 6'h2b : T388;
  assign T388 = T410 ? 6'h2c : T389;
  assign T389 = T409 ? 6'h2d : T390;
  assign T390 = T408 ? 6'h2e : T391;
  assign T391 = T407 ? 6'h2f : T392;
  assign T392 = T406 ? 6'h30 : T393;
  assign T393 = T405 ? 6'h31 : T394;
  assign T394 = T395 ? 6'h32 : 6'h33;
  assign T395 = T12[50];
  assign T12 = {T50, T13};
  assign T13 = {T25, T14};
  assign T14 = {T21, T15};
  assign T15 = {T20, T16};
  assign T16 = T17[1];
  assign T17 = T18[3:2];
  assign T18 = T19[19:16];
  assign T19 = T7[51:32];
  assign T20 = T17[0];
  assign T21 = {T24, T22};
  assign T22 = T23[1];
  assign T23 = T18[1:0];
  assign T24 = T23[0];
  assign T25 = T48 | T26;
  assign T26 = T27 & 16'haaaa;
  assign T27 = T28 << 1'h1;
  assign T28 = T29[14:0];
  assign T29 = T46 | T30;
  assign T30 = T31 & 16'hcccc;
  assign T31 = T32 << 2'h2;
  assign T32 = T33[13:0];
  assign T33 = T44 | T34;
  assign T34 = T35 & 16'hf0f0;
  assign T35 = T36 << 3'h4;
  assign T36 = T37[11:0];
  assign T37 = T42 | T38;
  assign T38 = T39 & 16'hff00;
  assign T39 = T40 << 4'h8;
  assign T40 = T41[7:0];
  assign T41 = T19[15:0];
  assign T42 = T396 & 16'hff;
  assign T396 = {8'h0, T43};
  assign T43 = T41 >> 4'h8;
  assign T44 = T397 & 16'hf0f;
  assign T397 = {4'h0, T45};
  assign T45 = T37 >> 3'h4;
  assign T46 = T398 & 16'h3333;
  assign T398 = {2'h0, T47};
  assign T47 = T33 >> 2'h2;
  assign T48 = T399 & 16'h5555;
  assign T399 = {1'h0, T49};
  assign T49 = T29 >> 1'h1;
  assign T50 = T79 | T51;
  assign T51 = T52 & 32'haaaaaaaa;
  assign T52 = T53 << 1'h1;
  assign T53 = T54[30:0];
  assign T54 = T77 | T55;
  assign T55 = T56 & 32'hcccccccc;
  assign T56 = T57 << 2'h2;
  assign T57 = T58[29:0];
  assign T58 = T75 | T59;
  assign T59 = T60 & 32'hf0f0f0f0;
  assign T60 = T61 << 3'h4;
  assign T61 = T62[27:0];
  assign T62 = T73 | T63;
  assign T63 = T64 & 32'hff00ff00;
  assign T64 = T65 << 4'h8;
  assign T65 = T66[23:0];
  assign T66 = T71 | T67;
  assign T67 = T68 & 32'hffff0000;
  assign T68 = T69 << 5'h10;
  assign T69 = T70[15:0];
  assign T70 = T7[31:0];
  assign T71 = T400 & 32'hffff;
  assign T400 = {16'h0, T72};
  assign T72 = T70 >> 5'h10;
  assign T73 = T401 & 32'hff00ff;
  assign T401 = {8'h0, T74};
  assign T74 = T66 >> 4'h8;
  assign T75 = T402 & 32'hf0f0f0f;
  assign T402 = {4'h0, T76};
  assign T76 = T62 >> 3'h4;
  assign T77 = T403 & 32'h33333333;
  assign T403 = {2'h0, T78};
  assign T78 = T58 >> 2'h2;
  assign T79 = T404 & 32'h55555555;
  assign T404 = {1'h0, T80};
  assign T80 = T54 >> 1'h1;
  assign T405 = T12[49];
  assign T406 = T12[48];
  assign T407 = T12[47];
  assign T408 = T12[46];
  assign T409 = T12[45];
  assign T410 = T12[44];
  assign T411 = T12[43];
  assign T412 = T12[42];
  assign T413 = T12[41];
  assign T414 = T12[40];
  assign T415 = T12[39];
  assign T416 = T12[38];
  assign T417 = T12[37];
  assign T418 = T12[36];
  assign T419 = T12[35];
  assign T420 = T12[34];
  assign T421 = T12[33];
  assign T422 = T12[32];
  assign T423 = T12[31];
  assign T424 = T12[30];
  assign T425 = T12[29];
  assign T426 = T12[28];
  assign T427 = T12[27];
  assign T428 = T12[26];
  assign T429 = T12[25];
  assign T430 = T12[24];
  assign T431 = T12[23];
  assign T432 = T12[22];
  assign T433 = T12[21];
  assign T434 = T12[20];
  assign T435 = T12[19];
  assign T436 = T12[18];
  assign T437 = T12[17];
  assign T438 = T12[16];
  assign T439 = T12[15];
  assign T440 = T12[14];
  assign T441 = T12[13];
  assign T442 = T12[12];
  assign T443 = T12[11];
  assign T444 = T12[10];
  assign T445 = T12[9];
  assign T446 = T12[8];
  assign T447 = T12[7];
  assign T448 = T12[6];
  assign T449 = T12[5];
  assign T450 = T12[4];
  assign T451 = T12[3];
  assign T452 = T12[2];
  assign T453 = T12[1];
  assign T454 = T12[0];
  assign T81 = T82 == 11'h0;
  assign T82 = io_b[62:52];
  assign T83 = T84 ^ 1'h1;
  assign T84 = T81 & T85;
  assign T85 = T7 == 52'h0;
  assign T86 = T87[8:0];
  assign T87 = T88;
  assign T88 = T89;
  assign T89 = {1'h0, T90};
  assign T90 = T91;
  assign T91 = T94 + T455;
  assign T455 = {1'h0, T92};
  assign T92 = 11'h400 | T456;
  assign T456 = {9'h0, T93};
  assign T93 = T81 ? 2'h2 : 2'h1;
  assign T94 = T81 ? T95 : T457;
  assign T457 = {1'h0, T82};
  assign T95 = T458 ^ 12'hfff;
  assign T458 = {6'h0, T344};
  assign T96 = {T106, T97};
  assign T97 = T103 | T459;
  assign T459 = {2'h0, T98};
  assign T98 = T99;
  assign T99 = T101 & T100;
  assign T100 = T85 ^ 1'h1;
  assign T101 = T102 == 2'h3;
  assign T102 = T91[11:10];
  assign T103 = T105 ? 3'h0 : T104;
  assign T104 = T87[11:9];
  assign T105 = T84;
  assign T106 = T107;
  assign T107 = io_b[63];
  assign T108 = {T204, T109};
  assign T109 = {T194, T110};
  assign T110 = T111[51:0];
  assign T111 = T112;
  assign T112 = {1'h0, T113};
  assign T113 = {T191, T114};
  assign T114 = T189 ? T116 : T115;
  assign T115 = io_a[51:0];
  assign T116 = T117 << 1'h1;
  assign T117 = T118[50:0];
  assign T118 = T115 << T460;
  assign T460 = T570 ? 1'h0 : T461;
  assign T461 = T569 ? 1'h1 : T462;
  assign T462 = T568 ? 2'h2 : T463;
  assign T463 = T567 ? 2'h3 : T464;
  assign T464 = T566 ? 3'h4 : T465;
  assign T465 = T565 ? 3'h5 : T466;
  assign T466 = T564 ? 3'h6 : T467;
  assign T467 = T563 ? 3'h7 : T468;
  assign T468 = T562 ? 4'h8 : T469;
  assign T469 = T561 ? 4'h9 : T470;
  assign T470 = T560 ? 4'ha : T471;
  assign T471 = T559 ? 4'hb : T472;
  assign T472 = T558 ? 4'hc : T473;
  assign T473 = T557 ? 4'hd : T474;
  assign T474 = T556 ? 4'he : T475;
  assign T475 = T555 ? 4'hf : T476;
  assign T476 = T554 ? 5'h10 : T477;
  assign T477 = T553 ? 5'h11 : T478;
  assign T478 = T552 ? 5'h12 : T479;
  assign T479 = T551 ? 5'h13 : T480;
  assign T480 = T550 ? 5'h14 : T481;
  assign T481 = T549 ? 5'h15 : T482;
  assign T482 = T548 ? 5'h16 : T483;
  assign T483 = T547 ? 5'h17 : T484;
  assign T484 = T546 ? 5'h18 : T485;
  assign T485 = T545 ? 5'h19 : T486;
  assign T486 = T544 ? 5'h1a : T487;
  assign T487 = T543 ? 5'h1b : T488;
  assign T488 = T542 ? 5'h1c : T489;
  assign T489 = T541 ? 5'h1d : T490;
  assign T490 = T540 ? 5'h1e : T491;
  assign T491 = T539 ? 5'h1f : T492;
  assign T492 = T538 ? 6'h20 : T493;
  assign T493 = T537 ? 6'h21 : T494;
  assign T494 = T536 ? 6'h22 : T495;
  assign T495 = T535 ? 6'h23 : T496;
  assign T496 = T534 ? 6'h24 : T497;
  assign T497 = T533 ? 6'h25 : T498;
  assign T498 = T532 ? 6'h26 : T499;
  assign T499 = T531 ? 6'h27 : T500;
  assign T500 = T530 ? 6'h28 : T501;
  assign T501 = T529 ? 6'h29 : T502;
  assign T502 = T528 ? 6'h2a : T503;
  assign T503 = T527 ? 6'h2b : T504;
  assign T504 = T526 ? 6'h2c : T505;
  assign T505 = T525 ? 6'h2d : T506;
  assign T506 = T524 ? 6'h2e : T507;
  assign T507 = T523 ? 6'h2f : T508;
  assign T508 = T522 ? 6'h30 : T509;
  assign T509 = T521 ? 6'h31 : T510;
  assign T510 = T511 ? 6'h32 : 6'h33;
  assign T511 = T120[50];
  assign T120 = {T158, T121};
  assign T121 = {T133, T122};
  assign T122 = {T129, T123};
  assign T123 = {T128, T124};
  assign T124 = T125[1];
  assign T125 = T126[3:2];
  assign T126 = T127[19:16];
  assign T127 = T115[51:32];
  assign T128 = T125[0];
  assign T129 = {T132, T130};
  assign T130 = T131[1];
  assign T131 = T126[1:0];
  assign T132 = T131[0];
  assign T133 = T156 | T134;
  assign T134 = T135 & 16'haaaa;
  assign T135 = T136 << 1'h1;
  assign T136 = T137[14:0];
  assign T137 = T154 | T138;
  assign T138 = T139 & 16'hcccc;
  assign T139 = T140 << 2'h2;
  assign T140 = T141[13:0];
  assign T141 = T152 | T142;
  assign T142 = T143 & 16'hf0f0;
  assign T143 = T144 << 3'h4;
  assign T144 = T145[11:0];
  assign T145 = T150 | T146;
  assign T146 = T147 & 16'hff00;
  assign T147 = T148 << 4'h8;
  assign T148 = T149[7:0];
  assign T149 = T127[15:0];
  assign T150 = T512 & 16'hff;
  assign T512 = {8'h0, T151};
  assign T151 = T149 >> 4'h8;
  assign T152 = T513 & 16'hf0f;
  assign T513 = {4'h0, T153};
  assign T153 = T145 >> 3'h4;
  assign T154 = T514 & 16'h3333;
  assign T514 = {2'h0, T155};
  assign T155 = T141 >> 2'h2;
  assign T156 = T515 & 16'h5555;
  assign T515 = {1'h0, T157};
  assign T157 = T137 >> 1'h1;
  assign T158 = T187 | T159;
  assign T159 = T160 & 32'haaaaaaaa;
  assign T160 = T161 << 1'h1;
  assign T161 = T162[30:0];
  assign T162 = T185 | T163;
  assign T163 = T164 & 32'hcccccccc;
  assign T164 = T165 << 2'h2;
  assign T165 = T166[29:0];
  assign T166 = T183 | T167;
  assign T167 = T168 & 32'hf0f0f0f0;
  assign T168 = T169 << 3'h4;
  assign T169 = T170[27:0];
  assign T170 = T181 | T171;
  assign T171 = T172 & 32'hff00ff00;
  assign T172 = T173 << 4'h8;
  assign T173 = T174[23:0];
  assign T174 = T179 | T175;
  assign T175 = T176 & 32'hffff0000;
  assign T176 = T177 << 5'h10;
  assign T177 = T178[15:0];
  assign T178 = T115[31:0];
  assign T179 = T516 & 32'hffff;
  assign T516 = {16'h0, T180};
  assign T180 = T178 >> 5'h10;
  assign T181 = T517 & 32'hff00ff;
  assign T517 = {8'h0, T182};
  assign T182 = T174 >> 4'h8;
  assign T183 = T518 & 32'hf0f0f0f;
  assign T518 = {4'h0, T184};
  assign T184 = T170 >> 3'h4;
  assign T185 = T519 & 32'h33333333;
  assign T519 = {2'h0, T186};
  assign T186 = T166 >> 2'h2;
  assign T187 = T520 & 32'h55555555;
  assign T520 = {1'h0, T188};
  assign T188 = T162 >> 1'h1;
  assign T521 = T120[49];
  assign T522 = T120[48];
  assign T523 = T120[47];
  assign T524 = T120[46];
  assign T525 = T120[45];
  assign T526 = T120[44];
  assign T527 = T120[43];
  assign T528 = T120[42];
  assign T529 = T120[41];
  assign T530 = T120[40];
  assign T531 = T120[39];
  assign T532 = T120[38];
  assign T533 = T120[37];
  assign T534 = T120[36];
  assign T535 = T120[35];
  assign T536 = T120[34];
  assign T537 = T120[33];
  assign T538 = T120[32];
  assign T539 = T120[31];
  assign T540 = T120[30];
  assign T541 = T120[29];
  assign T542 = T120[28];
  assign T543 = T120[27];
  assign T544 = T120[26];
  assign T545 = T120[25];
  assign T546 = T120[24];
  assign T547 = T120[23];
  assign T548 = T120[22];
  assign T549 = T120[21];
  assign T550 = T120[20];
  assign T551 = T120[19];
  assign T552 = T120[18];
  assign T553 = T120[17];
  assign T554 = T120[16];
  assign T555 = T120[15];
  assign T556 = T120[14];
  assign T557 = T120[13];
  assign T558 = T120[12];
  assign T559 = T120[11];
  assign T560 = T120[10];
  assign T561 = T120[9];
  assign T562 = T120[8];
  assign T563 = T120[7];
  assign T564 = T120[6];
  assign T565 = T120[5];
  assign T566 = T120[4];
  assign T567 = T120[3];
  assign T568 = T120[2];
  assign T569 = T120[1];
  assign T570 = T120[0];
  assign T189 = T190 == 11'h0;
  assign T190 = io_a[62:52];
  assign T191 = T192 ^ 1'h1;
  assign T192 = T189 & T193;
  assign T193 = T115 == 52'h0;
  assign T194 = T195[8:0];
  assign T195 = T196;
  assign T196 = T197;
  assign T197 = {1'h0, T198};
  assign T198 = T199;
  assign T199 = T202 + T571;
  assign T571 = {1'h0, T200};
  assign T200 = 11'h400 | T572;
  assign T572 = {9'h0, T201};
  assign T201 = T189 ? 2'h2 : 2'h1;
  assign T202 = T189 ? T203 : T573;
  assign T573 = {1'h0, T190};
  assign T203 = T574 ^ 12'hfff;
  assign T574 = {6'h0, T460};
  assign T204 = {T214, T205};
  assign T205 = T211 | T575;
  assign T575 = {2'h0, T206};
  assign T206 = T207;
  assign T207 = T209 & T208;
  assign T208 = T193 ^ 1'h1;
  assign T209 = T210 == 2'h3;
  assign T210 = T199[11:10];
  assign T211 = T213 ? 3'h0 : T212;
  assign T212 = T195[11:9];
  assign T213 = T192;
  assign T214 = T215;
  assign T215 = io_a[63];
  assign io_pass = T216;
  assign T216 = T218 & T217;
  assign T217 = io_actual_exceptionFlags == io_expected_exceptionFlags;
  assign T218 = T231 ? T226 : T219;
  assign T219 = T224 ? T221 : T220;
  assign T220 = io_actual_out == io_expected_recOut;
  assign T221 = T223 == T222;
  assign T222 = io_expected_recOut[64:61];
  assign T223 = io_actual_out[64:61];
  assign T224 = T225 == 3'h6;
  assign T225 = T223[2:0];
  assign T226 = T230 & T227;
  assign T227 = T229 == T228;
  assign T228 = io_expected_recOut[51:0];
  assign T229 = io_actual_out[51:0];
  assign T230 = T223 == T222;
  assign T231 = T234 | T232;
  assign T232 = T233 == 3'h7;
  assign T233 = T223[2:0];
  assign T234 = T235 == 3'h0;
  assign T235 = T223[2:0];
  assign io_check = 1'h1;
  assign io_actual_exceptionFlags = mulAddRecFN_io_exceptionFlags;
  assign io_actual_out = mulAddRecFN_io_out;
  assign io_expected_recOut = T236;
  assign T236 = {T332, T237};
  assign T237 = {T322, T238};
  assign T238 = T239[51:0];
  assign T239 = T240;
  assign T240 = {1'h0, T241};
  assign T241 = {T319, T242};
  assign T242 = T317 ? T244 : T243;
  assign T243 = io_expected_out[51:0];
  assign T244 = T245 << 1'h1;
  assign T245 = T246[50:0];
  assign T246 = T243 << T576;
  assign T576 = T686 ? 1'h0 : T577;
  assign T577 = T685 ? 1'h1 : T578;
  assign T578 = T684 ? 2'h2 : T579;
  assign T579 = T683 ? 2'h3 : T580;
  assign T580 = T682 ? 3'h4 : T581;
  assign T581 = T681 ? 3'h5 : T582;
  assign T582 = T680 ? 3'h6 : T583;
  assign T583 = T679 ? 3'h7 : T584;
  assign T584 = T678 ? 4'h8 : T585;
  assign T585 = T677 ? 4'h9 : T586;
  assign T586 = T676 ? 4'ha : T587;
  assign T587 = T675 ? 4'hb : T588;
  assign T588 = T674 ? 4'hc : T589;
  assign T589 = T673 ? 4'hd : T590;
  assign T590 = T672 ? 4'he : T591;
  assign T591 = T671 ? 4'hf : T592;
  assign T592 = T670 ? 5'h10 : T593;
  assign T593 = T669 ? 5'h11 : T594;
  assign T594 = T668 ? 5'h12 : T595;
  assign T595 = T667 ? 5'h13 : T596;
  assign T596 = T666 ? 5'h14 : T597;
  assign T597 = T665 ? 5'h15 : T598;
  assign T598 = T664 ? 5'h16 : T599;
  assign T599 = T663 ? 5'h17 : T600;
  assign T600 = T662 ? 5'h18 : T601;
  assign T601 = T661 ? 5'h19 : T602;
  assign T602 = T660 ? 5'h1a : T603;
  assign T603 = T659 ? 5'h1b : T604;
  assign T604 = T658 ? 5'h1c : T605;
  assign T605 = T657 ? 5'h1d : T606;
  assign T606 = T656 ? 5'h1e : T607;
  assign T607 = T655 ? 5'h1f : T608;
  assign T608 = T654 ? 6'h20 : T609;
  assign T609 = T653 ? 6'h21 : T610;
  assign T610 = T652 ? 6'h22 : T611;
  assign T611 = T651 ? 6'h23 : T612;
  assign T612 = T650 ? 6'h24 : T613;
  assign T613 = T649 ? 6'h25 : T614;
  assign T614 = T648 ? 6'h26 : T615;
  assign T615 = T647 ? 6'h27 : T616;
  assign T616 = T646 ? 6'h28 : T617;
  assign T617 = T645 ? 6'h29 : T618;
  assign T618 = T644 ? 6'h2a : T619;
  assign T619 = T643 ? 6'h2b : T620;
  assign T620 = T642 ? 6'h2c : T621;
  assign T621 = T641 ? 6'h2d : T622;
  assign T622 = T640 ? 6'h2e : T623;
  assign T623 = T639 ? 6'h2f : T624;
  assign T624 = T638 ? 6'h30 : T625;
  assign T625 = T637 ? 6'h31 : T626;
  assign T626 = T627 ? 6'h32 : 6'h33;
  assign T627 = T248[50];
  assign T248 = {T286, T249};
  assign T249 = {T261, T250};
  assign T250 = {T257, T251};
  assign T251 = {T256, T252};
  assign T252 = T253[1];
  assign T253 = T254[3:2];
  assign T254 = T255[19:16];
  assign T255 = T243[51:32];
  assign T256 = T253[0];
  assign T257 = {T260, T258};
  assign T258 = T259[1];
  assign T259 = T254[1:0];
  assign T260 = T259[0];
  assign T261 = T284 | T262;
  assign T262 = T263 & 16'haaaa;
  assign T263 = T264 << 1'h1;
  assign T264 = T265[14:0];
  assign T265 = T282 | T266;
  assign T266 = T267 & 16'hcccc;
  assign T267 = T268 << 2'h2;
  assign T268 = T269[13:0];
  assign T269 = T280 | T270;
  assign T270 = T271 & 16'hf0f0;
  assign T271 = T272 << 3'h4;
  assign T272 = T273[11:0];
  assign T273 = T278 | T274;
  assign T274 = T275 & 16'hff00;
  assign T275 = T276 << 4'h8;
  assign T276 = T277[7:0];
  assign T277 = T255[15:0];
  assign T278 = T628 & 16'hff;
  assign T628 = {8'h0, T279};
  assign T279 = T277 >> 4'h8;
  assign T280 = T629 & 16'hf0f;
  assign T629 = {4'h0, T281};
  assign T281 = T273 >> 3'h4;
  assign T282 = T630 & 16'h3333;
  assign T630 = {2'h0, T283};
  assign T283 = T269 >> 2'h2;
  assign T284 = T631 & 16'h5555;
  assign T631 = {1'h0, T285};
  assign T285 = T265 >> 1'h1;
  assign T286 = T315 | T287;
  assign T287 = T288 & 32'haaaaaaaa;
  assign T288 = T289 << 1'h1;
  assign T289 = T290[30:0];
  assign T290 = T313 | T291;
  assign T291 = T292 & 32'hcccccccc;
  assign T292 = T293 << 2'h2;
  assign T293 = T294[29:0];
  assign T294 = T311 | T295;
  assign T295 = T296 & 32'hf0f0f0f0;
  assign T296 = T297 << 3'h4;
  assign T297 = T298[27:0];
  assign T298 = T309 | T299;
  assign T299 = T300 & 32'hff00ff00;
  assign T300 = T301 << 4'h8;
  assign T301 = T302[23:0];
  assign T302 = T307 | T303;
  assign T303 = T304 & 32'hffff0000;
  assign T304 = T305 << 5'h10;
  assign T305 = T306[15:0];
  assign T306 = T243[31:0];
  assign T307 = T632 & 32'hffff;
  assign T632 = {16'h0, T308};
  assign T308 = T306 >> 5'h10;
  assign T309 = T633 & 32'hff00ff;
  assign T633 = {8'h0, T310};
  assign T310 = T302 >> 4'h8;
  assign T311 = T634 & 32'hf0f0f0f;
  assign T634 = {4'h0, T312};
  assign T312 = T298 >> 3'h4;
  assign T313 = T635 & 32'h33333333;
  assign T635 = {2'h0, T314};
  assign T314 = T294 >> 2'h2;
  assign T315 = T636 & 32'h55555555;
  assign T636 = {1'h0, T316};
  assign T316 = T290 >> 1'h1;
  assign T637 = T248[49];
  assign T638 = T248[48];
  assign T639 = T248[47];
  assign T640 = T248[46];
  assign T641 = T248[45];
  assign T642 = T248[44];
  assign T643 = T248[43];
  assign T644 = T248[42];
  assign T645 = T248[41];
  assign T646 = T248[40];
  assign T647 = T248[39];
  assign T648 = T248[38];
  assign T649 = T248[37];
  assign T650 = T248[36];
  assign T651 = T248[35];
  assign T652 = T248[34];
  assign T653 = T248[33];
  assign T654 = T248[32];
  assign T655 = T248[31];
  assign T656 = T248[30];
  assign T657 = T248[29];
  assign T658 = T248[28];
  assign T659 = T248[27];
  assign T660 = T248[26];
  assign T661 = T248[25];
  assign T662 = T248[24];
  assign T663 = T248[23];
  assign T664 = T248[22];
  assign T665 = T248[21];
  assign T666 = T248[20];
  assign T667 = T248[19];
  assign T668 = T248[18];
  assign T669 = T248[17];
  assign T670 = T248[16];
  assign T671 = T248[15];
  assign T672 = T248[14];
  assign T673 = T248[13];
  assign T674 = T248[12];
  assign T675 = T248[11];
  assign T676 = T248[10];
  assign T677 = T248[9];
  assign T678 = T248[8];
  assign T679 = T248[7];
  assign T680 = T248[6];
  assign T681 = T248[5];
  assign T682 = T248[4];
  assign T683 = T248[3];
  assign T684 = T248[2];
  assign T685 = T248[1];
  assign T686 = T248[0];
  assign T317 = T318 == 11'h0;
  assign T318 = io_expected_out[62:52];
  assign T319 = T320 ^ 1'h1;
  assign T320 = T317 & T321;
  assign T321 = T243 == 52'h0;
  assign T322 = T323[8:0];
  assign T323 = T324;
  assign T324 = T325;
  assign T325 = {1'h0, T326};
  assign T326 = T327;
  assign T327 = T330 + T687;
  assign T687 = {1'h0, T328};
  assign T328 = 11'h400 | T688;
  assign T688 = {9'h0, T329};
  assign T329 = T317 ? 2'h2 : 2'h1;
  assign T330 = T317 ? T331 : T689;
  assign T689 = {1'h0, T318};
  assign T331 = T690 ^ 12'hfff;
  assign T690 = {6'h0, T576};
  assign T332 = {T342, T333};
  assign T333 = T339 | T691;
  assign T691 = {2'h0, T334};
  assign T334 = T335;
  assign T335 = T337 & T336;
  assign T336 = T321 ^ 1'h1;
  assign T337 = T338 == 2'h3;
  assign T338 = T327[11:10];
  assign T339 = T341 ? 3'h0 : T340;
  assign T340 = T323[11:9];
  assign T341 = T320;
  assign T342 = T343;
  assign T343 = io_expected_out[63];
  MulAddRecFN mulAddRecFN(
       .io_op( 2'h0 ),
       .io_a( T108 ),
       .io_b( 65'h8000000000000000 ),
       .io_c( T0 ),
       .io_roundingMode( io_roundingMode ),
       .io_detectTininess( io_detectTininess ),
       .io_out( mulAddRecFN_io_out ),
       .io_exceptionFlags( mulAddRecFN_io_exceptionFlags )
  );
endmodule

